i_BEQ_0: assume property (i0[14:12] == 3'b000);
i_BEQ_1: assume property (i0[6:0] == 7'b1100011);
