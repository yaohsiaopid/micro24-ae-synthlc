i_ORI_0: assume property (i0[14:12] == 3'b110);
i_ORI_1: assume property (i0[11:7] != 5'd0);
i_ORI_2: assume property (i0[6:0] == 7'b0010011);
