i_BLT_0: assume property (i0[14:12] == 3'b100);
i_BLT_1: assume property (i0[6:0] == 7'b1100011);
