i_MULW_0: assume property (i0[31:25] == 7'b0000001);
i_MULW_1: assume property (i0[14:12] == 3'b000);
i_MULW_2: assume property (i0[11:7] != 5'd0);
i_MULW_3: assume property (i0[6:0] == 7'b0111011);
