i_BGE_0: assume property (i0[14:12] == 3'b101);
i_BGE_1: assume property (i0[6:0] == 7'b1100011);
