i_LHU_0: assume property (i0[14:12] == 3'b101);
i_LHU_1: assume property (i0[11:7] != 5'd0);
i_LHU_2: assume property (i0[6:0] == 7'b0000011);
