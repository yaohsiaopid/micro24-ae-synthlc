i_SH_0: assume property (i0[14:12] == 3'b001);
i_SH_1: assume property (i0[6:0] == 7'b0100011);
