`define SYSINSN
i_CSRRS_0: assume property (i0[14:12] == 3'b010);
i_CSRRS_2: assume property (i0[6:0] == 7'b1110011);
