i_ADDIW_0: assume property (i0[14:12] == 3'b000);
i_ADDIW_1: assume property (i0[11:7] != 5'd0);
i_ADDIW_2: assume property (i0[6:0] == 7'b0011011);
