group_0_i0: assume property (
(i0[11:7] != 5'd0 && i0[6:0] == 7'b1101111 &&  1'b1 ) || 
1'b0);
// 15||JAL
