i_SB_0: assume property (i0[14:12] == 3'b000);
i_SB_1: assume property (i0[6:0] == 7'b0100011);
