i_SRLI_0: assume property (i0[31:26] == 6'b000000);
i_SRLI_1: assume property (i0[14:12] == 3'b101);
i_SRLI_2: assume property (i0[11:7] != 5'd0);
i_SRLI_3: assume property (i0[6:0] == 7'b0010011);
