i_LH_0: assume property (i0[14:12] == 3'b001);
i_LH_1: assume property (i0[11:7] != 5'd0);
i_LH_2: assume property (i0[6:0] == 7'b0000011);
