i_SLLW_0: assume property (i0[31:25] == 7'b0000000);
i_SLLW_1: assume property (i0[14:12] == 3'b001);
i_SLLW_2: assume property (i0[11:7] != 5'd0);
i_SLLW_3: assume property (i0[6:0] == 7'b0111011);
