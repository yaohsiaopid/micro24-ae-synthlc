i_XORI_0: assume property (i0[14:12] == 3'b100);
i_XORI_1: assume property (i0[11:7] != 5'd0);
i_XORI_2: assume property (i0[6:0] == 7'b0010011);
