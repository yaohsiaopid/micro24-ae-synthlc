`define SYSINSN
i_CSRRSI_0: assume property (i0[14:12] == 3'b110);
i_CSRRSI_2: assume property (i0[6:0] == 7'b1110011);
