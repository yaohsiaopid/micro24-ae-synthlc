i_REMUW_0: assume property (i0[31:25] == 7'b0000001);
i_REMUW_1: assume property (i0[14:12] == 3'b111);
i_REMUW_2: assume property (i0[11:7] != 5'd0);
i_REMUW_3: assume property (i0[6:0] == 7'b0111011);
