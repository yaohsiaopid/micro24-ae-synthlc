i_SD_0: assume property (i0[14:12] == 3'b011);
i_SD_1: assume property (i0[6:0] == 7'b0100011);
