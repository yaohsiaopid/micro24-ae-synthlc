i_SLLI_0: assume property (i0[31:26] == 6'b000000);
i_SLLI_1: assume property (i0[14:12] == 3'b001);
i_SLLI_2: assume property (i0[11:7] != 5'd0);
i_SLLI_3: assume property (i0[6:0] == 7'b0010011);
