group_13_i0: assume property (
(i0[31:20] == 12'b000000000001 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[31:20] == 12'b000000000000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
1'b0);
// 13||EBREAK,ECALL
