group_10_i0: assume property (
(i0[14:12] == 3'b000 && i0[6:0] == 7'b1100111 &&  1'b1 ) || 
1'b0);
// JALR
