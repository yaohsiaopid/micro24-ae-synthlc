i_SRLW_0: assume property (i0[31:25] == 7'b0000000);
i_SRLW_1: assume property (i0[14:12] == 3'b101);
i_SRLW_2: assume property (i0[11:7] != 5'd0);
i_SRLW_3: assume property (i0[6:0] == 7'b0111011);
