group_2_i0: assume property (
((i0[31:25] == 7'b0000000) && (i0[14:12] == 3'b000) && (i0[11:7] != 5'd0) && (i0[6:0] == 7'b0110011) && 1'b1) || 
1'b0);
// ADD
