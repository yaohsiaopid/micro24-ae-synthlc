group_18_i0: assume property (
(i0[14:12] == 3'b000 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b001 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b010 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b100 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
(i0[14:12] == 3'b011 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0000011 &&  1'b1 ) || 
1'b0);
// LB,LH,LW,LBU,LHU,LWU,LD
