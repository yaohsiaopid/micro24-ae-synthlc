i_SRA_0: assume property (i0[31:25] == 7'b0100000);
i_SRA_1: assume property (i0[14:12] == 3'b101);
i_SRA_2: assume property (i0[11:7] != 5'd0);
i_SRA_3: assume property (i0[6:0] == 7'b0110011);
