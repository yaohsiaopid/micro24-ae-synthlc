i_BNE_0: assume property (i0[14:12] == 3'b001);
i_BNE_1: assume property (i0[6:0] == 7'b1100011);
