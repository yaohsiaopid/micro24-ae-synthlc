group_2_i0: assume property (
(i0[14:12] == 3'b000 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0011011 &&  1'b1 ) || 
(i0[31:25] == 7'b0000000 && i0[14:12] == 3'b001 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0011011 &&  1'b1 ) || 
(i0[31:25] == 7'b0000000 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0011011 &&  1'b1 ) || 
(i0[31:25] == 7'b0100000 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0011011 &&  1'b1 ) || 
1'b0);
// ADDIW,SLLIW,SRLIW,SRAIW
