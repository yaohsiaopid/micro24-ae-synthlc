group_8_i0: assume property (
(i0[14:12] == 3'b000 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[14:12] == 3'b010 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[14:12] == 3'b011 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[14:12] == 3'b100 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[14:12] == 3'b111 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[31:26] == 6'b000000 && i0[14:12] == 3'b001 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[31:26] == 6'b000000 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
(i0[31:26] == 6'b010000 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0010011 &&  1'b1 ) || 
1'b0);
// ADDI,SLTI,SLTIU,XORI,ORI,ANDI,SLLI,SRLI,SRAI
