i_JAL_0: assume property (i0[11:7] != 5'd0);
i_JAL_1: assume property (i0[6:0] == 7'b1101111);
