i_BLTU_0: assume property (i0[14:12] == 3'b110);
i_BLTU_1: assume property (i0[6:0] == 7'b1100011);
