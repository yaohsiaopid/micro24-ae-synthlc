i_AUIPC_0: assume property (i0[11:7] != 5'd0);
i_AUIPC_1: assume property (i0[6:0] == 7'b0010111);
