i_SLT_0: assume property (i0[31:25] == 7'b0000000);
i_SLT_1: assume property (i0[14:12] == 3'b010);
i_SLT_2: assume property (i0[11:7] != 5'd0);
i_SLT_3: assume property (i0[6:0] == 7'b0110011);
