i_LB_0: assume property (i0[14:12] == 3'b000);
i_LB_1: assume property (i0[11:7] != 5'd0);
i_LB_2: assume property (i0[6:0] == 7'b0000011);
