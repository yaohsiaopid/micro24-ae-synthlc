`define SYSINSN
i_CSRRWI_0: assume property (i0[14:12] == 3'b101);
i_CSRRWI_2: assume property (i0[6:0] == 7'b1110011);
