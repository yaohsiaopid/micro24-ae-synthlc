group_13_i0: assume property (
(i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[14:12] == 3'b111 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
1'b0);
