i_SRAI_0: assume property (i0[31:26] == 6'b010000);
i_SRAI_1: assume property (i0[14:12] == 3'b101);
i_SRAI_2: assume property (i0[11:7] != 5'd0);
i_SRAI_3: assume property (i0[6:0] == 7'b0010011);
