`define SYSINSN
i_CSRRC_0: assume property (i0[14:12] == 3'b011);
i_CSRRC_2: assume property (i0[6:0] == 7'b1110011);
