`define SYSINSN
i_CSRRW_0: assume property (i0[14:12] == 3'b001);
i_CSRRW_2: assume property (i0[6:0] == 7'b1110011);
