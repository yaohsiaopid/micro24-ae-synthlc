i_JALR_0: assume property (i0[14:12] == 3'b000);
i_JALR_1: assume property (i0[6:0] == 7'b1100111);
