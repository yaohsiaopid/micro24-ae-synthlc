i_MULHU_0: assume property (i0[31:25] == 7'b0000001);
i_MULHU_1: assume property (i0[14:12] == 3'b011);
i_MULHU_2: assume property (i0[11:7] != 5'd0);
i_MULHU_3: assume property (i0[6:0] == 7'b0110011);
