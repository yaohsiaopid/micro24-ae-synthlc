i_MULH_0: assume property (i0[31:25] == 7'b0000001);
i_MULH_1: assume property (i0[14:12] == 3'b001);
i_MULH_2: assume property (i0[11:7] != 5'd0);
i_MULH_3: assume property (i0[6:0] == 7'b0110011);
