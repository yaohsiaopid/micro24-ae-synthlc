group_4_i0: assume property (
((i0[14:12] == 3'b010) && (i0[6:0] == 7'b0100011) && 1'b1) ||
1'b0);
// SW
