i_BGEU_0: assume property (i0[14:12] == 3'b111);
i_BGEU_1: assume property (i0[6:0] == 7'b1100011);
