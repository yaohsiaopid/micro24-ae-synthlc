i_LUI_0: assume property (i0[11:7] != 5'd0);
i_LUI_1: assume property (i0[6:0] == 7'b0110111);
