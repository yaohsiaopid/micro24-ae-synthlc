group_0_i0: assume property (
(i0[31:20] == 12'b000000000001 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[11:7] != 5'd0 && i0[6:0] == 7'b0110111 &&  1'b1 ) || 
(i0[31:28] == 4'b0000 && i0[27:24] == 4'b0000 && i0[23:20] == 4'b0000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b001 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b0001111 &&  1'b1 ) || 
(i0[31:20] == 12'b000000000000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[11:7] != 5'd0 && i0[6:0] == 7'b1101111 &&  1'b1 ) || 
(i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[14:12] == 3'b111 && i0[11:7] != 5'd0 && i0[6:0] == 7'b1110011 &&  1'b1 ) || 
(i0[31:28] == 4'b0000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b0001111 &&  1'b1 ) || 
(i0[11:7] != 5'd0 && i0[6:0] == 7'b0010111 &&  1'b1 ) || 
1'b0);
// EBREAK,LUI,FENCEI,ECALL,JAL,CSRRSI,CSRRWI,CSRRCI,FENCE,AUIPC
