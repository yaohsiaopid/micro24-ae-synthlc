group_0_i0: assume property (
(i0[11:7] != 5'd0 && i0[6:0] == 7'b0110111 &&  1'b1 ) || 
(i0[11:7] != 5'd0 && i0[6:0] == 7'b0010111 &&  1'b1 ) || 
1'b0);
// 16||LUI,AUIPC
