group_11_i0: assume property (
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b100 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0111011 &&  1'b1 ) || // DIVW,      
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0111011 &&  1'b1 ) || // DIVUW,     
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0111011 &&  1'b1 ) || // REMW,      
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b110 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0110011 &&  1'b1 ) || // REM,       
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b111 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0110011 &&  1'b1 ) || // REMU,      
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b101 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0110011 &&  1'b1 ) || // DIVU,      
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b100 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0110011 &&  1'b1 ) || // DIV,       
    (i0[31:25] == 7'b0000001 && i0[14:12] == 3'b111 && i0[11:7] != 5'd0 && i0[6:0] == 7'b0111011 &&  1'b1 ) || // REMUW      
1'b0);
// DIV,DIVU,DIVUW,DIVW,REM,REMU,REMUW,REMW
