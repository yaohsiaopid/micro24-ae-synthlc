i_SUB_0: assume property (i0[31:25] == 7'b0100000);
i_SUB_1: assume property (i0[14:12] == 3'b000);
i_SUB_2: assume property (i0[11:7] != 5'd0);
i_SUB_3: assume property (i0[6:0] == 7'b0110011);
