module ariane(input clk_i
, input rst_ni
);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire _4776_;
  wire _4777_;
  wire _4778_;
  wire _4779_;
  wire _4780_;
  wire _4781_;
  wire _4782_;
  wire _4783_;
  wire _4784_;
  wire _4785_;
  wire _4786_;
  wire _4787_;
  wire _4788_;
  wire _4789_;
  wire _4790_;
  wire _4791_;
  wire _4792_;
  wire _4793_;
  wire _4794_;
  wire _4795_;
  wire _4796_;
  wire _4797_;
  wire _4798_;
  wire _4799_;
  wire _4800_;
  wire _4801_;
  wire _4802_;
  wire _4803_;
  wire _4804_;
  wire _4805_;
  wire _4806_;
  wire _4807_;
  wire _4808_;
  wire _4809_;
  wire _4810_;
  wire _4811_;
  wire _4812_;
  wire _4813_;
  wire _4814_;
  wire _4815_;
  wire _4816_;
  wire _4817_;
  wire _4818_;
  wire _4819_;
  wire _4820_;
  wire _4821_;
  wire _4822_;
  wire _4823_;
  wire _4824_;
  wire _4825_;
  wire _4826_;
  wire _4827_;
  wire _4828_;
  wire _4829_;
  wire _4830_;
  wire _4831_;
  wire _4832_;
  wire _4833_;
  wire _4834_;
  wire _4835_;
  wire _4836_;
  wire _4837_;
  wire _4838_;
  wire _4839_;
  wire _4840_;
  wire _4841_;
  wire _4842_;
  wire _4843_;
  wire _4844_;
  wire _4845_;
  wire _4846_;
  wire _4847_;
  wire _4848_;
  wire _4849_;
  wire _4850_;
  wire _4851_;
  wire _4852_;
  wire _4853_;
  wire _4854_;
  wire _4855_;
  wire _4856_;
  wire _4857_;
  wire _4858_;
  wire _4859_;
  wire _4860_;
  wire _4861_;
  wire _4862_;
  wire _4863_;
  wire _4864_;
  wire _4865_;
  wire _4866_;
  wire _4867_;
  wire _4868_;
  wire _4869_;
  wire _4870_;
  wire _4871_;
  wire _4872_;
  wire _4873_;
  wire _4874_;
  wire _4875_;
  wire _4876_;
  wire _4877_;
  wire _4878_;
  wire _4879_;
  wire _4880_;
  wire _4881_;
  wire _4882_;
  wire _4883_;
  wire _4884_;
  wire _4885_;
  wire _4886_;
  wire _4887_;
  wire _4888_;
  wire _4889_;
  wire _4890_;
  wire _4891_;
  wire _4892_;
  wire _4893_;
  wire _4894_;
  wire _4895_;
  wire _4896_;
  wire _4897_;
  wire _4898_;
  wire _4899_;
  wire _4900_;
  wire _4901_;
  wire _4902_;
  wire _4903_;
  wire _4904_;
  wire _4905_;
  wire _4906_;
  wire _4907_;
  wire _4908_;
  wire _4909_;
  wire _4910_;
  wire _4911_;
  wire _4912_;
  wire _4913_;
  wire _4914_;
  wire _4915_;
  wire _4916_;
  wire _4917_;
  wire _4918_;
  wire _4919_;
  wire _4920_;
  wire _4921_;
  wire _4922_;
  wire _4923_;
  wire _4924_;
  wire _4925_;
  wire _4926_;
  wire _4927_;
  wire _4928_;
  wire _4929_;
  wire _4930_;
  wire _4931_;
  wire _4932_;
  wire _4933_;
  wire _4934_;
  wire _4935_;
  wire _4936_;
  wire _4937_;
  wire _4938_;
  wire _4939_;
  wire _4940_;
  wire _4941_;
  wire _4942_;
  wire _4943_;
  wire _4944_;
  wire _4945_;
  wire _4946_;
  wire _4947_;
  wire _4948_;
  wire _4949_;
  wire _4950_;
  wire _4951_;
  wire _4952_;
  wire _4953_;
  wire _4954_;
  wire _4955_;
  wire _4956_;
  wire _4957_;
  wire _4958_;
  wire _4959_;
  wire _4960_;
  wire _4961_;
  wire _4962_;
  wire _4963_;
  wire _4964_;
  wire _4965_;
  wire _4966_;
  wire _4967_;
  wire _4968_;
  wire _4969_;
  wire _4970_;
  wire _4971_;
  wire _4972_;
  wire _4973_;
  wire _4974_;
  wire _4975_;
  wire _4976_;
  wire _4977_;
  wire _4978_;
  wire _4979_;
  wire _4980_;
  wire _4981_;
  wire _4982_;
  wire _4983_;
  wire _4984_;
  wire _4985_;
  wire _4986_;
  wire _4987_;
  wire _4988_;
  wire _4989_;
  wire _4990_;
  wire _4991_;
  wire _4992_;
  wire _4993_;
  wire _4994_;
  wire _4995_;
  wire _4996_;
  wire _4997_;
  wire _4998_;
  wire _4999_;
  wire _5000_;
  wire _5001_;
  wire _5002_;
  wire _5003_;
  wire _5004_;
  wire _5005_;
  wire _5006_;
  wire _5007_;
  wire _5008_;
  wire _5009_;
  wire _5010_;
  wire _5011_;
  wire _5012_;
  wire _5013_;
  wire _5014_;
  wire _5015_;
  wire _5016_;
  wire _5017_;
  wire _5018_;
  wire _5019_;
  wire _5020_;
  wire _5021_;
  wire _5022_;
  wire _5023_;
  wire _5024_;
  wire _5025_;
  wire _5026_;
  wire _5027_;
  wire _5028_;
  wire _5029_;
  wire _5030_;
  wire _5031_;
  wire _5032_;
  wire _5033_;
  wire _5034_;
  wire _5035_;
  wire _5036_;
  wire _5037_;
  wire _5038_;
  wire _5039_;
  wire _5040_;
  wire _5041_;
  wire _5042_;
  wire _5043_;
  wire _5044_;
  wire _5045_;
  wire _5046_;
  wire _5047_;
  wire _5048_;
  wire _5049_;
  wire _5050_;
  wire _5051_;
  wire _5052_;
  wire _5053_;
  wire _5054_;
  wire _5055_;
  wire _5056_;
  wire _5057_;
  wire _5058_;
  wire _5059_;
  wire _5060_;
  wire _5061_;
  wire _5062_;
  wire _5063_;
  wire _5064_;
  wire _5065_;
  wire _5066_;
  wire _5067_;
  wire _5068_;
  wire _5069_;
  wire _5070_;
  wire _5071_;
  wire _5072_;
  wire _5073_;
  wire _5074_;
  wire _5075_;
  wire _5076_;
  wire _5077_;
  wire _5078_;
  wire _5079_;
  wire _5080_;
  wire _5081_;
  wire _5082_;
  wire _5083_;
  wire _5084_;
  wire _5085_;
  wire _5086_;
  wire _5087_;
  wire _5088_;
  wire _5089_;
  wire _5090_;
  wire _5091_;
  wire _5092_;
  wire _5093_;
  wire _5094_;
  wire _5095_;
  wire _5096_;
  wire _5097_;
  wire _5098_;
  wire _5099_;
  wire _5100_;
  wire _5101_;
  wire _5102_;
  wire _5103_;
  wire _5104_;
  wire _5105_;
  wire _5106_;
  wire _5107_;
  wire _5108_;
  wire _5109_;
  wire _5110_;
  wire _5111_;
  wire _5112_;
  wire _5113_;
  wire _5114_;
  wire _5115_;
  wire _5116_;
  wire _5117_;
  wire _5118_;
  wire _5119_;
  wire _5120_;
  wire _5121_;
  wire _5122_;
  wire _5123_;
  wire _5124_;
  wire _5125_;
  wire _5126_;
  wire _5127_;
  wire _5128_;
  wire _5129_;
  wire _5130_;
  wire _5131_;
  wire _5132_;
  wire _5133_;
  wire _5134_;
  wire _5135_;
  wire _5136_;
  wire _5137_;
  wire _5138_;
  wire _5139_;
  wire _5140_;
  wire _5141_;
  wire _5142_;
  wire _5143_;
  wire _5144_;
  wire _5145_;
  wire _5146_;
  wire _5147_;
  wire _5148_;
  wire _5149_;
  wire _5150_;
  wire _5151_;
  wire _5152_;
  wire _5153_;
  wire _5154_;
  wire _5155_;
  wire _5156_;
  wire _5157_;
  wire _5158_;
  wire _5159_;
  wire _5160_;
  wire _5161_;
  wire _5162_;
  wire _5163_;
  wire _5164_;
  wire _5165_;
  wire _5166_;
  wire _5167_;
  wire _5168_;
  wire _5169_;
  wire _5170_;
  wire _5171_;
  wire _5172_;
  wire _5173_;
  wire _5174_;
  wire _5175_;
  wire _5176_;
  wire _5177_;
  wire _5178_;
  wire _5179_;
  wire _5180_;
  wire _5181_;
  wire _5182_;
  wire _5183_;
  wire _5184_;
  wire _5185_;
  wire _5186_;
  wire _5187_;
  wire _5188_;
  wire _5189_;
  wire _5190_;
  wire _5191_;
  wire _5192_;
  wire _5193_;
  wire _5194_;
  wire _5195_;
  wire _5196_;
  wire _5197_;
  wire _5198_;
  wire _5199_;
  wire _5200_;
  wire _5201_;
  wire _5202_;
  wire _5203_;
  wire _5204_;
  wire _5205_;
  wire _5206_;
  wire _5207_;
  wire _5208_;
  wire _5209_;
  wire _5210_;
  wire _5211_;
  wire _5212_;
  wire _5213_;
  wire _5214_;
  wire _5215_;
  wire _5216_;
  wire _5217_;
  wire _5218_;
  wire _5219_;
  wire _5220_;
  wire _5221_;
  wire _5222_;
  wire _5223_;
  wire _5224_;
  wire _5225_;
  wire _5226_;
  wire _5227_;
  wire _5228_;
  wire _5229_;
  wire _5230_;
  wire _5231_;
  wire _5232_;
  wire _5233_;
  wire _5234_;
  wire _5235_;
  wire _5236_;
  wire _5237_;
  wire _5238_;
  wire _5239_;
  wire _5240_;
  wire _5241_;
  wire _5242_;
  wire _5243_;
  wire _5244_;
  wire _5245_;
  wire _5246_;
  wire _5247_;
  wire _5248_;
  wire _5249_;
  wire _5250_;
  wire _5251_;
  wire _5252_;
  wire _5253_;
  wire _5254_;
  wire _5255_;
  wire _5256_;
  wire _5257_;
  wire _5258_;
  wire _5259_;
  wire _5260_;
  wire _5261_;
  wire _5262_;
  wire _5263_;
  wire _5264_;
  wire _5265_;
  wire _5266_;
  wire _5267_;
  wire _5268_;
  wire _5269_;
  wire _5270_;
  wire _5271_;
  wire _5272_;
  wire _5273_;
  wire _5274_;
  wire _5275_;
  wire _5276_;
  wire _5277_;
  wire _5278_;
  wire _5279_;
  wire _5280_;
  wire _5281_;
  wire _5282_;
  wire _5283_;
  wire _5284_;
  wire _5285_;
  wire _5286_;
  wire _5287_;
  wire _5288_;
  wire _5289_;
  wire _5290_;
  wire _5291_;
  wire _5292_;
  wire _5293_;
  wire _5294_;
  wire _5295_;
  wire _5296_;
  wire _5297_;
  wire _5298_;
  wire _5299_;
  wire _5300_;
  wire _5301_;
  wire _5302_;
  wire _5303_;
  wire _5304_;
  wire _5305_;
  wire _5306_;
  wire _5307_;
  wire _5308_;
  wire _5309_;
  wire _5310_;
  wire _5311_;
  wire _5312_;
  wire _5313_;
  wire _5314_;
  wire _5315_;
  wire _5316_;
  wire _5317_;
  wire _5318_;
  wire _5319_;
  wire _5320_;
  wire _5321_;
  wire _5322_;
  wire _5323_;
  wire _5324_;
  wire _5325_;
  wire _5326_;
  wire _5327_;
  wire _5328_;
  wire _5329_;
  wire _5330_;
  wire _5331_;
  wire _5332_;
  wire _5333_;
  wire _5334_;
  wire _5335_;
  wire _5336_;
  wire _5337_;
  wire _5338_;
  wire _5339_;
  wire _5340_;
  wire _5341_;
  wire _5342_;
  wire _5343_;
  wire _5344_;
  wire _5345_;
  wire _5346_;
  wire _5347_;
  wire _5348_;
  wire _5349_;
  wire _5350_;
  wire _5351_;
  wire _5352_;
  wire _5353_;
  wire _5354_;
  wire _5355_;
  wire _5356_;
  wire _5357_;
  wire _5358_;
  wire _5359_;
  wire _5360_;
  wire _5361_;
  wire _5362_;
  wire _5363_;
  wire _5364_;
  wire _5365_;
  wire _5366_;
  wire _5367_;
  wire _5368_;
  wire _5369_;
  wire _5370_;
  wire _5371_;
  wire _5372_;
  wire _5373_;
  wire _5374_;
  wire _5375_;
  wire _5376_;
  wire _5377_;
  wire _5378_;
  wire _5379_;
  wire _5380_;
  wire _5381_;
  wire _5382_;
  wire _5383_;
  wire _5384_;
  wire _5385_;
  wire _5386_;
  wire _5387_;
  wire _5388_;
  wire _5389_;
  wire _5390_;
  wire _5391_;
  wire _5392_;
  wire _5393_;
  wire _5394_;
  wire _5395_;
  wire _5396_;
  wire _5397_;
  wire _5398_;
  wire _5399_;
  wire _5400_;
  wire _5401_;
  wire _5402_;
  wire _5403_;
  wire _5404_;
  wire _5405_;
  wire _5406_;
  wire _5407_;
  wire _5408_;
  wire _5409_;
  wire _5410_;
  wire _5411_;
  wire _5412_;
  wire _5413_;
  wire _5414_;
  wire _5415_;
  wire _5416_;
  wire _5417_;
  wire _5418_;
  wire _5419_;
  wire _5420_;
  wire _5421_;
  wire _5422_;
  wire _5423_;
  wire _5424_;
  wire _5425_;
  wire _5426_;
  wire _5427_;
  wire _5428_;
  wire _5429_;
  wire _5430_;
  wire _5431_;
  wire _5432_;
  wire _5433_;
  wire _5434_;
  wire _5435_;
  wire _5436_;
  wire _5437_;
  wire _5438_;
  wire _5439_;
  wire _5440_;
  wire _5441_;
  wire _5442_;
  wire _5443_;
  wire _5444_;
  wire _5445_;
  wire _5446_;
  wire _5447_;
  wire _5448_;
  wire _5449_;
  wire _5450_;
  wire _5451_;
  wire _5452_;
  wire _5453_;
  wire _5454_;
  wire _5455_;
  wire _5456_;
  wire _5457_;
  wire _5458_;
  wire _5459_;
  wire _5460_;
  wire _5461_;
  wire _5462_;
  wire _5463_;
  wire _5464_;
  wire _5465_;
  wire _5466_;
  wire _5467_;
  wire _5468_;
  wire _5469_;
  wire _5470_;
  wire _5471_;
  wire _5472_;
  wire _5473_;
  wire _5474_;
  wire _5475_;
  wire _5476_;
  wire _5477_;
  wire _5478_;
  wire _5479_;
  wire _5480_;
  wire _5481_;
  wire _5482_;
  wire _5483_;
  wire _5484_;
  wire _5485_;
  wire _5486_;
  wire _5487_;
  wire _5488_;
  wire _5489_;
  wire _5490_;
  wire _5491_;
  wire _5492_;
  wire _5493_;
  wire _5494_;
  wire _5495_;
  wire _5496_;
  wire _5497_;
  wire _5498_;
  wire _5499_;
  wire _5500_;
  wire _5501_;
  wire _5502_;
  wire _5503_;
  wire _5504_;
  wire _5505_;
  wire _5506_;
  wire _5507_;
  wire _5508_;
  wire _5509_;
  wire _5510_;
  wire _5511_;
  wire _5512_;
  wire _5513_;
  wire _5514_;
  wire _5515_;
  wire _5516_;
  wire _5517_;
  wire _5518_;
  wire _5519_;
  wire _5520_;
  wire _5521_;
  wire _5522_;
  wire _5523_;
  wire _5524_;
  wire _5525_;
  wire _5526_;
  wire _5527_;
  wire _5528_;
  wire _5529_;
  wire _5530_;
  wire _5531_;
  wire _5532_;
  wire _5533_;
  wire _5534_;
  wire _5535_;
  wire _5536_;
  wire _5537_;
  wire _5538_;
  wire _5539_;
  wire _5540_;
  wire _5541_;
  wire _5542_;
  wire _5543_;
  wire _5544_;
  wire _5545_;
  wire _5546_;
  wire _5547_;
  wire _5548_;
  wire _5549_;
  wire _5550_;
  wire _5551_;
  wire _5552_;
  wire _5553_;
  wire _5554_;
  wire _5555_;
  wire _5556_;
  wire _5557_;
  wire _5558_;
  wire _5559_;
  wire _5560_;
  wire _5561_;
  wire _5562_;
  wire _5563_;
  wire _5564_;
  wire _5565_;
  wire _5566_;
  wire _5567_;
  wire _5568_;
  wire _5569_;
  wire _5570_;
  wire _5571_;
  wire _5572_;
  wire _5573_;
  wire _5574_;
  wire _5575_;
  wire _5576_;
  wire _5577_;
  wire _5578_;
  wire _5579_;
  wire _5580_;
  wire _5581_;
  wire _5582_;
  wire _5583_;
  wire _5584_;
  wire _5585_;
  wire _5586_;
  wire _5587_;
  wire _5588_;
  wire _5589_;
  wire _5590_;
  wire _5591_;
  wire _5592_;
  wire _5593_;
  wire _5594_;
  wire _5595_;
  wire _5596_;
  wire _5597_;
  wire _5598_;
  wire _5599_;
  wire _5600_;
  wire _5601_;
  wire _5602_;
  wire _5603_;
  wire _5604_;
  wire _5605_;
  wire _5606_;
  wire _5607_;
  wire _5608_;
  wire _5609_;
  wire _5610_;
  wire _5611_;
  wire _5612_;
  wire _5613_;
  wire _5614_;
  wire _5615_;
  wire _5616_;
  wire _5617_;
  wire _5618_;
  wire _5619_;
  wire _5620_;
  wire _5621_;
  wire _5622_;
  wire _5623_;
  wire _5624_;
  wire _5625_;
  wire _5626_;
  wire _5627_;
  wire _5628_;
  wire _5629_;
  wire _5630_;
  wire _5631_;
  wire _5632_;
  wire _5633_;
  wire _5634_;
  wire _5635_;
  wire _5636_;
  wire _5637_;
  wire _5638_;
  wire _5639_;
  wire _5640_;
  wire _5641_;
  wire _5642_;
  wire _5643_;
  wire _5644_;
  wire _5645_;
  wire _5646_;
  wire _5647_;
  wire _5648_;
  wire _5649_;
  wire _5650_;
  wire _5651_;
  wire _5652_;
  wire _5653_;
  wire _5654_;
  wire _5655_;
  wire _5656_;
  wire _5657_;
  wire _5658_;
  wire _5659_;
  wire _5660_;
  wire _5661_;
  wire _5662_;
  wire _5663_;
  wire _5664_;
  wire _5665_;
  wire _5666_;
  wire _5667_;
  wire _5668_;
  wire _5669_;
  wire _5670_;
  wire _5671_;
  wire _5672_;
  wire _5673_;
  wire _5674_;
  wire _5675_;
  wire _5676_;
  wire _5677_;
  wire _5678_;
  wire _5679_;
  wire _5680_;
  wire _5681_;
  wire _5682_;
  wire _5683_;
  wire _5684_;
  wire _5685_;
  wire _5686_;
  wire _5687_;
  wire _5688_;
  wire _5689_;
  wire _5690_;
  wire _5691_;
  wire _5692_;
  wire _5693_;
  wire _5694_;
  wire _5695_;
  wire _5696_;
  wire _5697_;
  wire _5698_;
  wire _5699_;
  wire _5700_;
  wire _5701_;
  wire _5702_;
  wire _5703_;
  wire _5704_;
  wire _5705_;
  wire _5706_;
  wire _5707_;
  wire _5708_;
  wire _5709_;
  wire _5710_;
  wire _5711_;
  wire _5712_;
  wire _5713_;
  wire _5714_;
  wire _5715_;
  wire _5716_;
  wire _5717_;
  wire _5718_;
  wire _5719_;
  wire _5720_;
  wire _5721_;
  wire _5722_;
  wire _5723_;
  wire _5724_;
  wire _5725_;
  wire _5726_;
  wire _5727_;
  wire _5728_;
  wire _5729_;
  wire _5730_;
  wire _5731_;
  wire _5732_;
  wire _5733_;
  wire _5734_;
  wire _5735_;
  wire _5736_;
  wire _5737_;
  wire _5738_;
  wire _5739_;
  wire _5740_;
  wire _5741_;
  wire _5742_;
  wire _5743_;
  wire _5744_;
  wire _5745_;
  wire _5746_;
  wire _5747_;
  wire _5748_;
  wire _5749_;
  wire _5750_;
  wire _5751_;
  wire _5752_;
  wire _5753_;
  wire _5754_;
  wire _5755_;
  wire _5756_;
  wire _5757_;
  wire _5758_;
  wire _5759_;
  wire _5760_;
  wire _5761_;
  wire _5762_;
  wire _5763_;
  wire _5764_;
  wire _5765_;
  wire _5766_;
  wire _5767_;
  wire _5768_;
  wire _5769_;
  wire _5770_;
  wire _5771_;
  wire _5772_;
  wire _5773_;
  wire _5774_;
  wire _5775_;
  wire _5776_;
  wire _5777_;
  wire _5778_;
  wire _5779_;
  wire _5780_;
  wire _5781_;
  wire _5782_;
  wire _5783_;
  wire _5784_;
  wire _5785_;
  wire _5786_;
  wire _5787_;
  wire _5788_;
  wire _5789_;
  wire _5790_;
  wire _5791_;
  wire _5792_;
  wire _5793_;
  wire _5794_;
  wire _5795_;
  wire _5796_;
  wire _5797_;
  wire _5798_;
  wire _5799_;
  wire _5800_;
  wire _5801_;
  wire _5802_;
  wire _5803_;
  wire _5804_;
  wire _5805_;
  wire _5806_;
  wire _5807_;
  wire _5808_;
  wire _5809_;
  wire _5810_;
  wire _5811_;
  wire _5812_;
  wire _5813_;
  wire _5814_;
  wire _5815_;
  wire _5816_;
  wire _5817_;
  wire _5818_;
  wire _5819_;
  wire _5820_;
  wire _5821_;
  wire _5822_;
  wire _5823_;
  wire _5824_;
  wire _5825_;
  wire _5826_;
  wire _5827_;
  wire _5828_;
  wire _5829_;
  wire _5830_;
  wire _5831_;
  wire _5832_;
  wire _5833_;
  wire _5834_;
  wire _5835_;
  wire _5836_;
  wire _5837_;
  wire _5838_;
  wire _5839_;
  wire _5840_;
  wire _5841_;
  wire _5842_;
  wire _5843_;
  wire _5844_;
  wire _5845_;
  wire _5846_;
  wire _5847_;
  wire _5848_;
  wire _5849_;
  wire _5850_;
  wire _5851_;
  wire _5852_;
  wire _5853_;
  wire _5854_;
  wire _5855_;
  wire _5856_;
  wire _5857_;
  wire _5858_;
  wire _5859_;
  wire _5860_;
  wire _5861_;
  wire _5862_;
  wire _5863_;
  wire _5864_;
  wire _5865_;
  wire _5866_;
  wire _5867_;
  wire _5868_;
  wire _5869_;
  wire _5870_;
  wire _5871_;
  wire _5872_;
  wire _5873_;
  wire _5874_;
  wire _5875_;
  wire _5876_;
  wire _5877_;
  wire _5878_;
  wire _5879_;
  wire _5880_;
  wire _5881_;
  wire _5882_;
  wire _5883_;
  wire _5884_;
  wire _5885_;
  wire _5886_;
  wire _5887_;
  wire _5888_;
  wire _5889_;
  wire _5890_;
  wire _5891_;
  wire _5892_;
  wire _5893_;
  wire _5894_;
  wire _5895_;
  wire _5896_;
  wire _5897_;
  wire _5898_;
  wire _5899_;
  wire _5900_;
  wire _5901_;
  wire _5902_;
  wire _5903_;
  wire _5904_;
  wire _5905_;
  wire _5906_;
  wire _5907_;
  wire _5908_;
  wire _5909_;
  wire _5910_;
  wire _5911_;
  wire _5912_;
  wire _5913_;
  wire _5914_;
  wire _5915_;
  wire _5916_;
  wire _5917_;
  wire _5918_;
  wire _5919_;
  wire _5920_;
  wire _5921_;
  wire _5922_;
  wire _5923_;
  wire _5924_;
  wire _5925_;
  wire _5926_;
  wire _5927_;
  wire _5928_;
  wire _5929_;
  wire _5930_;
  wire _5931_;
  wire _5932_;
  wire _5933_;
  wire _5934_;
  wire _5935_;
  wire _5936_;
  wire _5937_;
  wire _5938_;
  wire _5939_;
  wire _5940_;
  wire _5941_;
  wire _5942_;
  wire _5943_;
  wire _5944_;
  wire _5945_;
  wire _5946_;
  wire _5947_;
  wire _5948_;
  wire _5949_;
  wire _5950_;
  wire _5951_;
  wire _5952_;
  wire _5953_;
  wire _5954_;
  wire _5955_;
  wire _5956_;
  wire _5957_;
  wire _5958_;
  wire _5959_;
  wire _5960_;
  wire _5961_;
  wire _5962_;
  wire _5963_;
  wire _5964_;
  wire _5965_;
  wire _5966_;
  wire _5967_;
  wire _5968_;
  wire _5969_;
  wire _5970_;
  wire _5971_;
  wire _5972_;
  wire _5973_;
  wire _5974_;
  wire _5975_;
  wire _5976_;
  wire _5977_;
  wire _5978_;
  wire _5979_;
  wire _5980_;
  wire _5981_;
  wire _5982_;
  wire _5983_;
  wire _5984_;
  wire _5985_;
  wire _5986_;
  wire _5987_;
  wire _5988_;
  wire _5989_;
  wire _5990_;
  wire _5991_;
  wire _5992_;
  wire _5993_;
  wire _5994_;
  wire _5995_;
  wire _5996_;
  wire _5997_;
  wire _5998_;
  wire _5999_;
  wire _6000_;
  wire _6001_;
  wire _6002_;
  wire _6003_;
  wire _6004_;
  wire _6005_;
  wire _6006_;
  wire _6007_;
  wire _6008_;
  wire _6009_;
  wire _6010_;
  wire _6011_;
  wire _6012_;
  wire _6013_;
  wire _6014_;
  wire _6015_;
  wire _6016_;
  wire _6017_;
  wire _6018_;
  wire _6019_;
  wire _6020_;
  wire _6021_;
  wire _6022_;
  wire _6023_;
  wire _6024_;
  wire _6025_;
  wire _6026_;
  wire _6027_;
  wire _6028_;
  wire _6029_;
  wire _6030_;
  wire _6031_;
  wire _6032_;
  wire _6033_;
  wire _6034_;
  wire _6035_;
  wire _6036_;
  wire _6037_;
  wire _6038_;
  wire _6039_;
  wire _6040_;
  wire _6041_;
  wire _6042_;
  wire _6043_;
  wire _6044_;
  wire _6045_;
  wire _6046_;
  wire _6047_;
  wire _6048_;
  wire _6049_;
  wire _6050_;
  wire _6051_;
  wire _6052_;
  wire _6053_;
  wire _6054_;
  wire _6055_;
  wire _6056_;
  wire _6057_;
  wire _6058_;
  wire _6059_;
  wire _6060_;
  wire _6061_;
  wire _6062_;
  wire _6063_;
  wire _6064_;
  wire _6065_;
  wire _6066_;
  wire _6067_;
  wire _6068_;
  wire _6069_;
  wire _6070_;
  wire _6071_;
  wire _6072_;
  wire _6073_;
  wire _6074_;
  wire _6075_;
  wire _6076_;
  wire _6077_;
  wire _6078_;
  wire _6079_;
  wire _6080_;
  wire _6081_;
  wire _6082_;
  wire _6083_;
  wire _6084_;
  wire _6085_;
  wire _6086_;
  wire _6087_;
  wire _6088_;
  wire _6089_;
  wire _6090_;
  wire _6091_;
  wire _6092_;
  wire _6093_;
  wire _6094_;
  wire _6095_;
  wire _6096_;
  wire _6097_;
  wire _6098_;
  wire _6099_;
  wire _6100_;
  wire _6101_;
  wire _6102_;
  wire _6103_;
  wire _6104_;
  wire _6105_;
  wire _6106_;
  wire _6107_;
  wire _6108_;
  wire _6109_;
  wire _6110_;
  wire _6111_;
  wire _6112_;
  wire _6113_;
  wire _6114_;
  wire _6115_;
  wire _6116_;
  wire _6117_;
  wire _6118_;
  wire _6119_;
  wire _6120_;
  wire _6121_;
  wire _6122_;
  wire _6123_;
  wire _6124_;
  wire _6125_;
  wire _6126_;
  wire _6127_;
  wire _6128_;
  wire _6129_;
  wire _6130_;
  wire _6131_;
  wire _6132_;
  wire _6133_;
  wire _6134_;
  wire _6135_;
  wire _6136_;
  wire _6137_;
  wire _6138_;
  wire _6139_;
  wire _6140_;
  wire _6141_;
  wire _6142_;
  wire _6143_;
  wire _6144_;
  wire _6145_;
  wire _6146_;
  wire _6147_;
  wire _6148_;
  wire _6149_;
  wire _6150_;
  wire _6151_;
  wire _6152_;
  wire _6153_;
  wire _6154_;
  wire _6155_;
  wire _6156_;
  wire _6157_;
  wire _6158_;
  wire _6159_;
  wire _6160_;
  wire _6161_;
  wire _6162_;
  wire _6163_;
  wire _6164_;
  wire _6165_;
  wire _6166_;
  wire _6167_;
  wire _6168_;
  wire _6169_;
  wire _6170_;
  wire _6171_;
  wire _6172_;
  wire _6173_;
  wire _6174_;
  wire _6175_;
  wire _6176_;
  wire _6177_;
  wire _6178_;
  wire _6179_;
  wire _6180_;
  wire _6181_;
  wire _6182_;
  wire _6183_;
  wire _6184_;
  wire _6185_;
  wire _6186_;
  wire _6187_;
  wire _6188_;
  wire _6189_;
  wire _6190_;
  wire _6191_;
  wire _6192_;
  wire _6193_;
  wire _6194_;
  wire _6195_;
  wire _6196_;
  wire _6197_;
  wire _6198_;
  wire _6199_;
  wire _6200_;
  wire _6201_;
  wire _6202_;
  wire _6203_;
  wire _6204_;
  wire _6205_;
  wire _6206_;
  wire _6207_;
  wire _6208_;
  wire _6209_;
  wire _6210_;
  wire _6211_;
  wire _6212_;
  wire _6213_;
  wire _6214_;
  wire _6215_;
  wire _6216_;
  wire _6217_;
  wire _6218_;
  wire _6219_;
  wire _6220_;
  wire _6221_;
  wire _6222_;
  wire _6223_;
  wire _6224_;
  wire _6225_;
  wire _6226_;
  wire _6227_;
  wire _6228_;
  wire _6229_;
  wire _6230_;
  wire _6231_;
  wire _6232_;
  wire _6233_;
  wire _6234_;
  wire _6235_;
  wire _6236_;
  wire _6237_;
  wire _6238_;
  wire _6239_;
  wire _6240_;
  wire _6241_;
  wire _6242_;
  wire _6243_;
  wire _6244_;
  wire _6245_;
  wire _6246_;
  wire _6247_;
  wire _6248_;
  wire _6249_;
  wire _6250_;
  wire _6251_;
  wire _6252_;
  wire _6253_;
  wire _6254_;
  wire _6255_;
  wire _6256_;
  wire _6257_;
  wire _6258_;
  wire _6259_;
  wire _6260_;
  wire _6261_;
  wire _6262_;
  wire _6263_;
  wire _6264_;
  wire _6265_;
  wire _6266_;
  wire _6267_;
  wire _6268_;
  wire _6269_;
  wire _6270_;
  wire _6271_;
  wire _6272_;
  wire _6273_;
  wire _6274_;
  wire _6275_;
  wire _6276_;
  wire _6277_;
  wire _6278_;
  wire _6279_;
  wire _6280_;
  wire _6281_;
  wire _6282_;
  wire _6283_;
  wire _6284_;
  wire _6285_;
  wire _6286_;
  wire _6287_;
  wire _6288_;
  wire _6289_;
  wire _6290_;
  wire _6291_;
  wire _6292_;
  wire _6293_;
  wire _6294_;
  wire _6295_;
  wire _6296_;
  wire _6297_;
  wire _6298_;
  wire _6299_;
  wire _6300_;
  wire _6301_;
  wire _6302_;
  wire _6303_;
  wire _6304_;
  wire _6305_;
  wire _6306_;
  wire _6307_;
  wire _6308_;
  wire _6309_;
  wire _6310_;
  wire _6311_;
  wire _6312_;
  wire _6313_;
  wire _6314_;
  wire _6315_;
  wire _6316_;
  wire _6317_;
  wire _6318_;
  wire _6319_;
  wire _6320_;
  wire _6321_;
  wire _6322_;
  wire _6323_;
  wire _6324_;
  wire _6325_;
  wire _6326_;
  wire _6327_;
  wire _6328_;
  wire _6329_;
  wire _6330_;
  wire _6331_;
  wire _6332_;
  wire _6333_;
  wire _6334_;
  wire _6335_;
  wire _6336_;
  wire _6337_;
  wire _6338_;
  wire _6339_;
  wire _6340_;
  wire _6341_;
  wire _6342_;
  wire _6343_;
  wire _6344_;
  wire _6345_;
  wire _6346_;
  wire _6347_;
  wire _6348_;
  wire _6349_;
  wire _6350_;
  wire _6351_;
  wire _6352_;
  wire _6353_;
  wire _6354_;
  wire _6355_;
  wire _6356_;
  wire _6357_;
  wire _6358_;
  wire _6359_;
  wire _6360_;
  wire _6361_;
  wire _6362_;
  wire _6363_;
  wire _6364_;
  wire _6365_;
  wire _6366_;
  wire _6367_;
  wire _6368_;
  wire _6369_;
  wire _6370_;
  wire _6371_;
  wire _6372_;
  wire _6373_;
  wire _6374_;
  wire _6375_;
  wire _6376_;
  wire _6377_;
  wire _6378_;
  wire _6379_;
  wire _6380_;
  wire _6381_;
  wire _6382_;
  wire _6383_;
  wire _6384_;
  wire _6385_;
  wire _6386_;
  wire _6387_;
  wire _6388_;
  wire _6389_;
  wire _6390_;
  wire _6391_;
  wire _6392_;
  wire _6393_;
  wire _6394_;
  wire _6395_;
  wire _6396_;
  wire _6397_;
  wire _6398_;
  wire _6399_;
  wire _6400_;
  wire _6401_;
  wire _6402_;
  wire _6403_;
  wire _6404_;
  wire _6405_;
  wire _6406_;
  wire _6407_;
  wire _6408_;
  wire _6409_;
  wire _6410_;
  wire _6411_;
  wire _6412_;
  wire _6413_;
  wire _6414_;
  wire _6415_;
  wire _6416_;
  wire _6417_;
  wire _6418_;
  wire _6419_;
  wire _6420_;
  wire _6421_;
  wire _6422_;
  wire _6423_;
  wire _6424_;
  wire _6425_;
  wire _6426_;
  wire _6427_;
  wire _6428_;
  wire _6429_;
  wire _6430_;
  wire _6431_;
  wire _6432_;
  wire _6433_;
  wire _6434_;
  wire _6435_;
  wire _6436_;
  wire _6437_;
  wire _6438_;
  wire _6439_;
  wire _6440_;
  wire _6441_;
  wire _6442_;
  wire _6443_;
  wire _6444_;
  wire _6445_;
  wire _6446_;
  wire _6447_;
  wire _6448_;
  wire _6449_;
  wire _6450_;
  wire _6451_;
  wire _6452_;
  wire _6453_;
  wire _6454_;
  wire _6455_;
  wire _6456_;
  wire _6457_;
  wire _6458_;
  wire _6459_;
  wire _6460_;
  wire _6461_;
  wire _6462_;
  wire _6463_;
  wire _6464_;
  wire _6465_;
  wire _6466_;
  wire _6467_;
  wire _6468_;
  wire _6469_;
  wire _6470_;
  wire _6471_;
  wire _6472_;
  wire _6473_;
  wire _6474_;
  wire _6475_;
  wire _6476_;
  wire _6477_;
  wire _6478_;
  wire _6479_;
  wire _6480_;
  wire _6481_;
  wire _6482_;
  wire _6483_;
  wire _6484_;
  wire _6485_;
  wire _6486_;
  wire _6487_;
  wire _6488_;
  wire _6489_;
  wire _6490_;
  wire _6491_;
  wire _6492_;
  wire _6493_;
  wire _6494_;
  wire _6495_;
  wire _6496_;
  wire _6497_;
  wire _6498_;
  wire _6499_;
  wire _6500_;
  wire _6501_;
  wire _6502_;
  wire _6503_;
  wire _6504_;
  wire _6505_;
  wire _6506_;
  wire _6507_;
  wire _6508_;
  wire _6509_;
  wire _6510_;
  wire _6511_;
  wire _6512_;
  wire _6513_;
  wire _6514_;
  wire _6515_;
  wire _6516_;
  wire _6517_;
  wire _6518_;
  wire _6519_;
  wire _6520_;
  wire _6521_;
  wire _6522_;
  wire _6523_;
  wire _6524_;
  wire _6525_;
  wire _6526_;
  wire _6527_;
  wire _6528_;
  wire _6529_;
  wire _6530_;
  wire _6531_;
  wire _6532_;
  wire _6533_;
  wire _6534_;
  wire _6535_;
  wire _6536_;
  wire _6537_;
  wire _6538_;
  wire _6539_;
  wire _6540_;
  wire _6541_;
  wire _6542_;
  wire _6543_;
  wire _6544_;
  wire _6545_;
  wire _6546_;
  wire _6547_;
  wire _6548_;
  wire _6549_;
  wire _6550_;
  wire _6551_;
  wire _6552_;
  wire _6553_;
  wire _6554_;
  wire _6555_;
  wire _6556_;
  wire _6557_;
  wire _6558_;
  wire _6559_;
  wire _6560_;
  wire _6561_;
  wire _6562_;
  wire _6563_;
  wire _6564_;
  wire _6565_;
  wire _6566_;
  wire _6567_;
  wire _6568_;
  wire _6569_;
  wire _6570_;
  wire _6571_;
  wire _6572_;
  wire _6573_;
  wire _6574_;
  wire _6575_;
  wire _6576_;
  wire _6577_;
  wire _6578_;
  wire _6579_;
  wire _6580_;
  wire _6581_;
  wire _6582_;
  wire _6583_;
  wire _6584_;
  wire _6585_;
  wire _6586_;
  wire _6587_;
  wire _6588_;
  wire _6589_;
  wire _6590_;
  wire _6591_;
  wire _6592_;
  wire _6593_;
  wire _6594_;
  wire _6595_;
  wire _6596_;
  wire _6597_;
  wire _6598_;
  wire _6599_;
  wire _6600_;
  wire _6601_;
  wire _6602_;
  wire _6603_;
  wire _6604_;
  wire _6605_;
  wire _6606_;
  wire _6607_;
  wire _6608_;
  wire _6609_;
  wire _6610_;
  wire _6611_;
  wire _6612_;
  wire _6613_;
  wire _6614_;
  wire _6615_;
  wire _6616_;
  wire _6617_;
  wire _6618_;
  wire _6619_;
  wire _6620_;
  wire _6621_;
  wire _6622_;
  wire _6623_;
  wire _6624_;
  wire _6625_;
  wire _6626_;
  wire _6627_;
  wire _6628_;
  wire _6629_;
  wire _6630_;
  wire _6631_;
  wire _6632_;
  wire _6633_;
  wire _6634_;
  wire _6635_;
  wire _6636_;
  wire _6637_;
  wire _6638_;
  wire _6639_;
  wire _6640_;
  wire _6641_;
  wire _6642_;
  wire _6643_;
  wire _6644_;
  wire _6645_;
  wire _6646_;
  wire _6647_;
  wire _6648_;
  wire _6649_;
  wire _6650_;
  wire _6651_;
  wire _6652_;
  wire _6653_;
  wire _6654_;
  wire _6655_;
  wire _6656_;
  wire _6657_;
  wire _6658_;
  wire _6659_;
  wire _6660_;
  wire _6661_;
  wire _6662_;
  wire _6663_;
  wire _6664_;
  wire _6665_;
  wire _6666_;
  wire _6667_;
  wire _6668_;
  wire _6669_;
  wire _6670_;
  wire _6671_;
  wire _6672_;
  wire _6673_;
  wire _6674_;
  wire _6675_;
  wire _6676_;
  wire _6677_;
  wire _6678_;
  wire _6679_;
  wire _6680_;
  wire _6681_;
  wire _6682_;
  wire _6683_;
  wire _6684_;
  wire _6685_;
  wire _6686_;
  wire _6687_;
  wire _6688_;
  wire _6689_;
  wire _6690_;
  wire _6691_;
  wire _6692_;
  wire _6693_;
  wire _6694_;
  wire _6695_;
  wire _6696_;
  wire _6697_;
  wire _6698_;
  wire _6699_;
  wire _6700_;
  wire _6701_;
  wire _6702_;
  wire _6703_;
  wire _6704_;
  wire _6705_;
  wire _6706_;
  wire _6707_;
  wire _6708_;
  wire _6709_;
  wire _6710_;
  wire _6711_;
  wire _6712_;
  wire _6713_;
  wire _6714_;
  wire _6715_;
  wire _6716_;
  wire _6717_;
  wire _6718_;
  wire _6719_;
  wire _6720_;
  wire _6721_;
  wire _6722_;
  wire _6723_;
  wire _6724_;
  wire _6725_;
  wire _6726_;
  wire _6727_;
  wire _6728_;
  wire _6729_;
  wire _6730_;
  wire _6731_;
  wire _6732_;
  wire _6733_;
  wire _6734_;
  wire _6735_;
  wire _6736_;
  wire _6737_;
  wire _6738_;
  wire _6739_;
  wire _6740_;
  wire _6741_;
  wire _6742_;
  wire _6743_;
  wire _6744_;
  wire _6745_;
  wire _6746_;
  wire _6747_;
  wire _6748_;
  wire _6749_;
  wire _6750_;
  wire _6751_;
  wire _6752_;
  wire _6753_;
  wire _6754_;
  wire _6755_;
  wire _6756_;
  wire _6757_;
  wire _6758_;
  wire _6759_;
  wire _6760_;
  wire _6761_;
  wire _6762_;
  wire _6763_;
  wire _6764_;
  wire _6765_;
  wire _6766_;
  wire _6767_;
  wire _6768_;
  wire _6769_;
  wire _6770_;
  wire _6771_;
  wire _6772_;
  wire _6773_;
  wire _6774_;
  wire _6775_;
  wire _6776_;
  wire _6777_;
  wire _6778_;
  wire _6779_;
  wire _6780_;
  wire _6781_;
  wire _6782_;
  wire _6783_;
  wire _6784_;
  wire _6785_;
  wire _6786_;
  wire _6787_;
  wire _6788_;
  wire _6789_;
  wire _6790_;
  wire _6791_;
  wire _6792_;
  wire _6793_;
  wire _6794_;
  wire _6795_;
  wire _6796_;
  wire _6797_;
  wire _6798_;
  wire _6799_;
  wire _6800_;
  wire _6801_;
  wire _6802_;
  wire _6803_;
  wire _6804_;
  wire _6805_;
  wire _6806_;
  wire _6807_;
  wire _6808_;
  wire _6809_;
  wire _6810_;
  wire _6811_;
  wire _6812_;
  wire _6813_;
  wire _6814_;
  wire _6815_;
  wire _6816_;
  wire _6817_;
  wire _6818_;
  wire _6819_;
  wire _6820_;
  wire _6821_;
  wire _6822_;
  wire _6823_;
  wire _6824_;
  wire _6825_;
  wire _6826_;
  wire _6827_;
  wire _6828_;
  wire _6829_;
  wire _6830_;
  wire _6831_;
  wire _6832_;
  wire _6833_;
  wire _6834_;
  wire _6835_;
  wire _6836_;
  wire _6837_;
  wire _6838_;
  wire _6839_;
  wire _6840_;
  wire _6841_;
  wire _6842_;
  wire _6843_;
  wire _6844_;
  wire _6845_;
  wire _6846_;
  wire _6847_;
  wire _6848_;
  wire _6849_;
  wire _6850_;
  wire _6851_;
  wire _6852_;
  wire _6853_;
  wire _6854_;
  wire _6855_;
  wire _6856_;
  wire _6857_;
  wire _6858_;
  wire _6859_;
  wire _6860_;
  wire _6861_;
  wire _6862_;
  wire _6863_;
  wire _6864_;
  wire _6865_;
  wire _6866_;
  wire _6867_;
  wire _6868_;
  wire _6869_;
  wire _6870_;
  wire _6871_;
  wire _6872_;
  wire _6873_;
  wire _6874_;
  wire _6875_;
  wire _6876_;
  wire _6877_;
  wire _6878_;
  wire _6879_;
  wire _6880_;
  wire _6881_;
  wire _6882_;
  wire _6883_;
  wire _6884_;
  wire _6885_;
  wire _6886_;
  wire _6887_;
  wire _6888_;
  wire _6889_;
  wire _6890_;
  wire _6891_;
  wire _6892_;
  wire _6893_;
  wire _6894_;
  wire _6895_;
  wire _6896_;
  wire _6897_;
  wire _6898_;
  wire _6899_;
  wire _6900_;
  wire _6901_;
  wire _6902_;
  wire _6903_;
  wire _6904_;
  wire _6905_;
  wire _6906_;
  wire _6907_;
  wire _6908_;
  wire _6909_;
  wire _6910_;
  wire _6911_;
  wire _6912_;
  wire _6913_;
  wire _6914_;
  wire _6915_;
  wire _6916_;
  wire _6917_;
  wire _6918_;
  wire _6919_;
  wire _6920_;
  wire _6921_;
  wire _6922_;
  wire _6923_;
  wire _6924_;
  wire _6925_;
  wire _6926_;
  wire _6927_;
  wire _6928_;
  wire _6929_;
  wire _6930_;
  wire _6931_;
  wire _6932_;
  wire _6933_;
  wire _6934_;
  wire _6935_;
  wire _6936_;
  wire _6937_;
  wire _6938_;
  wire _6939_;
  wire _6940_;
  wire _6941_;
  wire _6942_;
  wire _6943_;
  wire _6944_;
  wire _6945_;
  wire _6946_;
  wire _6947_;
  wire _6948_;
  wire _6949_;
  wire _6950_;
  wire _6951_;
  wire _6952_;
  wire _6953_;
  wire _6954_;
  wire _6955_;
  wire _6956_;
  wire _6957_;
  wire _6958_;
  wire _6959_;
  wire _6960_;
  wire _6961_;
  wire _6962_;
  wire _6963_;
  wire _6964_;
  wire _6965_;
  wire _6966_;
  wire _6967_;
  wire _6968_;
  wire _6969_;
  wire _6970_;
  wire _6971_;
  wire _6972_;
  wire _6973_;
  wire _6974_;
  wire _6975_;
  wire _6976_;
  wire _6977_;
  wire _6978_;
  wire _6979_;
  wire _6980_;
  wire _6981_;
  wire _6982_;
  wire _6983_;
  wire _6984_;
  wire _6985_;
  wire _6986_;
  wire _6987_;
  wire _6988_;
  wire _6989_;
  wire _6990_;
  wire _6991_;
  wire _6992_;
  wire _6993_;
  wire _6994_;
  wire _6995_;
  wire _6996_;
  wire _6997_;
  wire _6998_;
  wire _6999_;
  wire _7000_;
  wire _7001_;
  wire _7002_;
  wire _7003_;
  wire _7004_;
  wire _7005_;
  wire _7006_;
  wire _7007_;
  wire _7008_;
  wire _7009_;
  wire _7010_;
  wire _7011_;
  wire _7012_;
  wire _7013_;
  wire _7014_;
  wire _7015_;
  wire _7016_;
  wire _7017_;
  wire _7018_;
  wire _7019_;
  wire _7020_;
  wire _7021_;
  wire _7022_;
  wire _7023_;
  wire _7024_;
  wire _7025_;
  wire _7026_;
  wire _7027_;
  wire _7028_;
  wire _7029_;
  wire _7030_;
  wire _7031_;
  wire _7032_;
  wire _7033_;
  wire _7034_;
  wire _7035_;
  wire _7036_;
  wire _7037_;
  wire _7038_;
  wire _7039_;
  wire _7040_;
  wire _7041_;
  wire _7042_;
  wire _7043_;
  wire _7044_;
  wire _7045_;
  wire _7046_;
  wire _7047_;
  wire _7048_;
  wire _7049_;
  wire _7050_;
  wire _7051_;
  wire _7052_;
  wire _7053_;
  wire _7054_;
  wire _7055_;
  wire _7056_;
  wire _7057_;
  wire _7058_;
  wire _7059_;
  wire _7060_;
  wire _7061_;
  wire _7062_;
  wire _7063_;
  wire _7064_;
  wire _7065_;
  wire _7066_;
  wire _7067_;
  wire _7068_;
  wire _7069_;
  wire _7070_;
  wire _7071_;
  wire _7072_;
  wire _7073_;
  wire _7074_;
  wire _7075_;
  wire _7076_;
  wire _7077_;
  wire _7078_;
  wire _7079_;
  wire _7080_;
  wire _7081_;
  wire _7082_;
  wire _7083_;
  wire _7084_;
  wire _7085_;
  wire _7086_;
  wire _7087_;
  wire _7088_;
  wire _7089_;
  wire _7090_;
  wire _7091_;
  wire _7092_;
  wire _7093_;
  wire _7094_;
  wire _7095_;
  wire _7096_;
  wire _7097_;
  wire _7098_;
  wire _7099_;
  wire _7100_;
  wire _7101_;
  wire _7102_;
  wire _7103_;
  wire _7104_;
  wire _7105_;
  wire _7106_;
  wire _7107_;
  wire _7108_;
  wire _7109_;
  wire _7110_;
  wire _7111_;
  wire _7112_;
  wire _7113_;
  wire _7114_;
  wire _7115_;
  wire _7116_;
  wire _7117_;
  wire _7118_;
  wire _7119_;
  wire _7120_;
  wire _7121_;
  wire _7122_;
  wire _7123_;
  wire _7124_;
  wire _7125_;
  wire _7126_;
  wire _7127_;
  wire _7128_;
  wire _7129_;
  wire _7130_;
  wire _7131_;
  wire _7132_;
  wire _7133_;
  wire _7134_;
  wire _7135_;
  wire _7136_;
  wire _7137_;
  wire _7138_;
  wire _7139_;
  wire _7140_;
  wire _7141_;
  wire _7142_;
  wire _7143_;
  wire _7144_;
  wire _7145_;
  wire _7146_;
  wire _7147_;
  wire _7148_;
  wire _7149_;
  wire _7150_;
  wire _7151_;
  wire _7152_;
  wire _7153_;
  wire _7154_;
  wire _7155_;
  wire _7156_;
  wire _7157_;
  wire _7158_;
  wire _7159_;
  wire _7160_;
  wire _7161_;
  wire _7162_;
  wire _7163_;
  wire _7164_;
  wire _7165_;
  wire _7166_;
  wire _7167_;
  wire _7168_;
  wire _7169_;
  wire _7170_;
  wire _7171_;
  wire _7172_;
  wire _7173_;
  wire _7174_;
  wire _7175_;
  wire _7176_;
  wire _7177_;
  wire _7178_;
  wire _7179_;
  wire _7180_;
  wire _7181_;
  wire _7182_;
  wire _7183_;
  wire _7184_;
  wire _7185_;
  wire _7186_;
  wire _7187_;
  wire _7188_;
  wire _7189_;
  wire _7190_;
  wire _7191_;
  wire _7192_;
  wire _7193_;
  wire _7194_;
  wire _7195_;
  wire _7196_;
  wire _7197_;
  wire _7198_;
  wire _7199_;
  wire _7200_;
  wire _7201_;
  wire _7202_;
  wire _7203_;
  wire _7204_;
  wire _7205_;
  wire _7206_;
  wire _7207_;
  wire _7208_;
  wire _7209_;
  wire _7210_;
  wire _7211_;
  wire _7212_;
  wire _7213_;
  wire _7214_;
  wire _7215_;
  wire _7216_;
  wire _7217_;
  wire _7218_;
  wire _7219_;
  wire _7220_;
  wire _7221_;
  wire _7222_;
  wire _7223_;
  wire _7224_;
  wire _7225_;
  wire _7226_;
  wire _7227_;
  wire _7228_;
  wire _7229_;
  wire _7230_;
  wire _7231_;
  wire _7232_;
  wire _7233_;
  wire _7234_;
  wire _7235_;
  wire _7236_;
  wire _7237_;
  wire _7238_;
  wire _7239_;
  wire _7240_;
  wire _7241_;
  wire _7242_;
  wire _7243_;
  wire _7244_;
  wire _7245_;
  wire _7246_;
  wire _7247_;
  wire _7248_;
  wire _7249_;
  wire _7250_;
  wire _7251_;
  wire _7252_;
  wire _7253_;
  wire _7254_;
  wire _7255_;
  wire _7256_;
  wire _7257_;
  wire _7258_;
  wire _7259_;
  wire _7260_;
  wire _7261_;
  wire _7262_;
  wire _7263_;
  wire _7264_;
  wire _7265_;
  wire _7266_;
  wire _7267_;
  wire _7268_;
  wire _7269_;
  wire _7270_;
  wire _7271_;
  wire _7272_;
  wire _7273_;
  wire _7274_;
  wire _7275_;
  wire _7276_;
  wire _7277_;
  wire _7278_;
  wire _7279_;
  wire _7280_;
  wire _7281_;
  wire _7282_;
  wire _7283_;
  wire _7284_;
  wire _7285_;
  wire _7286_;
  wire _7287_;
  wire _7288_;
  wire _7289_;
  wire _7290_;
  wire _7291_;
  wire _7292_;
  wire _7293_;
  wire _7294_;
  wire _7295_;
  wire _7296_;
  wire _7297_;
  wire _7298_;
  wire _7299_;
  wire _7300_;
  wire _7301_;
  wire _7302_;
  wire _7303_;
  wire _7304_;
  wire _7305_;
  wire _7306_;
  wire _7307_;
  wire _7308_;
  wire _7309_;
  wire _7310_;
  wire _7311_;
  wire _7312_;
  wire _7313_;
  wire _7314_;
  wire _7315_;
  wire _7316_;
  wire _7317_;
  wire _7318_;
  wire _7319_;
  wire _7320_;
  wire _7321_;
  wire _7322_;
  wire _7323_;
  wire _7324_;
  wire _7325_;
  wire _7326_;
  wire _7327_;
  wire _7328_;
  wire _7329_;
  wire _7330_;
  wire _7331_;
  wire _7332_;
  wire _7333_;
  wire _7334_;
  wire _7335_;
  wire _7336_;
  wire _7337_;
  wire _7338_;
  wire _7339_;
  wire _7340_;
  wire _7341_;
  wire _7342_;
  wire _7343_;
  wire _7344_;
  wire _7345_;
  wire _7346_;
  wire _7347_;
  wire _7348_;
  wire _7349_;
  wire _7350_;
  wire _7351_;
  wire _7352_;
  wire _7353_;
  wire _7354_;
  wire _7355_;
  wire _7356_;
  wire _7357_;
  wire _7358_;
  wire _7359_;
  wire _7360_;
  wire _7361_;
  wire _7362_;
  wire _7363_;
  wire _7364_;
  wire _7365_;
  wire _7366_;
  wire _7367_;
  wire _7368_;
  wire _7369_;
  wire _7370_;
  wire _7371_;
  wire _7372_;
  wire _7373_;
  wire _7374_;
  wire _7375_;
  wire _7376_;
  wire _7377_;
  wire _7378_;
  wire _7379_;
  wire _7380_;
  wire _7381_;
  wire _7382_;
  wire _7383_;
  wire _7384_;
  wire _7385_;
  wire _7386_;
  wire _7387_;
  wire _7388_;
  wire _7389_;
  wire _7390_;
  wire _7391_;
  wire _7392_;
  wire _7393_;
  wire _7394_;
  wire _7395_;
  wire _7396_;
  wire _7397_;
  wire _7398_;
  wire _7399_;
  wire _7400_;
  wire _7401_;
  wire _7402_;
  wire _7403_;
  wire _7404_;
  wire _7405_;
  wire _7406_;
  wire _7407_;
  wire _7408_;
  wire _7409_;
  wire _7410_;
  wire _7411_;
  wire _7412_;
  wire _7413_;
  wire _7414_;
  wire _7415_;
  wire _7416_;
  wire _7417_;
  wire _7418_;
  wire _7419_;
  wire _7420_;
  wire _7421_;
  wire _7422_;
  wire _7423_;
  wire _7424_;
  wire _7425_;
  wire _7426_;
  wire _7427_;
  wire _7428_;
  wire _7429_;
  wire _7430_;
  wire _7431_;
  wire _7432_;
  wire _7433_;
  wire _7434_;
  wire _7435_;
  wire _7436_;
  wire _7437_;
  wire _7438_;
  wire _7439_;
  wire _7440_;
  wire _7441_;
  wire _7442_;
  wire _7443_;
  wire _7444_;
  wire _7445_;
  wire _7446_;
  wire _7447_;
  wire _7448_;
  wire _7449_;
  wire _7450_;
  wire _7451_;
  wire _7452_;
  wire _7453_;
  wire _7454_;
  wire _7455_;
  wire _7456_;
  wire _7457_;
  wire _7458_;
  wire _7459_;
  wire _7460_;
  wire _7461_;
  wire _7462_;
  wire _7463_;
  wire _7464_;
  wire _7465_;
  wire _7466_;
  wire _7467_;
  wire _7468_;
  wire _7469_;
  wire _7470_;
  wire _7471_;
  wire _7472_;
  wire _7473_;
  wire _7474_;
  wire _7475_;
  wire _7476_;
  wire _7477_;
  wire _7478_;
  wire _7479_;
  wire _7480_;
  wire _7481_;
  wire _7482_;
  wire _7483_;
  wire _7484_;
  wire _7485_;
  wire _7486_;
  wire _7487_;
  wire _7488_;
  wire _7489_;
  wire _7490_;
  wire _7491_;
  wire _7492_;
  wire _7493_;
  wire _7494_;
  wire _7495_;
  wire _7496_;
  wire _7497_;
  wire _7498_;
  wire _7499_;
  wire _7500_;
  wire _7501_;
  wire _7502_;
  wire _7503_;
  wire _7504_;
  wire _7505_;
  wire _7506_;
  wire _7507_;
  wire _7508_;
  wire _7509_;
  wire _7510_;
  wire _7511_;
  wire _7512_;
  wire _7513_;
  wire _7514_;
  wire _7515_;
  wire _7516_;
  wire _7517_;
  wire _7518_;
  wire _7519_;
  wire _7520_;
  wire _7521_;
  wire _7522_;
  wire _7523_;
  wire _7524_;
  wire _7525_;
  wire _7526_;
  wire _7527_;
  wire _7528_;
  wire _7529_;
  wire _7530_;
  wire _7531_;
  wire _7532_;
  wire _7533_;
  wire _7534_;
  wire _7535_;
  wire _7536_;
  wire _7537_;
  wire _7538_;
  wire _7539_;
  wire _7540_;
  wire _7541_;
  wire _7542_;
  wire _7543_;
  wire _7544_;
  wire _7545_;
  wire _7546_;
  wire _7547_;
  wire _7548_;
  wire _7549_;
  wire _7550_;
  wire _7551_;
  wire _7552_;
  wire _7553_;
  wire _7554_;
  wire _7555_;
  wire _7556_;
  wire _7557_;
  wire _7558_;
  wire _7559_;
  wire _7560_;
  wire _7561_;
  wire _7562_;
  wire _7563_;
  wire _7564_;
  wire _7565_;
  wire _7566_;
  wire _7567_;
  wire _7568_;
  wire _7569_;
  wire _7570_;
  wire _7571_;
  wire _7572_;
  wire _7573_;
  wire _7574_;
  wire _7575_;
  wire _7576_;
  wire _7577_;
  wire _7578_;
  wire _7579_;
  wire _7580_;
  wire _7581_;
  wire _7582_;
  wire _7583_;
  wire _7584_;
  wire _7585_;
  wire _7586_;
  wire _7587_;
  wire _7588_;
  wire _7589_;
  wire _7590_;
  wire _7591_;
  wire _7592_;
  wire _7593_;
  wire _7594_;
  wire _7595_;
  wire _7596_;
  wire _7597_;
  wire _7598_;
  wire _7599_;
  wire _7600_;
  wire _7601_;
  wire _7602_;
  wire _7603_;
  wire _7604_;
  wire _7605_;
  wire _7606_;
  wire _7607_;
  wire _7608_;
  wire _7609_;
  wire _7610_;
  wire _7611_;
  wire _7612_;
  wire _7613_;
  wire _7614_;
  wire _7615_;
  wire _7616_;
  wire _7617_;
  wire _7618_;
  wire _7619_;
  wire _7620_;
  wire _7621_;
  wire _7622_;
  wire _7623_;
  wire _7624_;
  wire _7625_;
  wire _7626_;
  wire _7627_;
  wire _7628_;
  wire _7629_;
  wire _7630_;
  wire _7631_;
  wire _7632_;
  wire _7633_;
  wire _7634_;
  wire _7635_;
  wire _7636_;
  wire _7637_;
  wire _7638_;
  wire _7639_;
  wire _7640_;
  wire _7641_;
  wire _7642_;
  wire _7643_;
  wire _7644_;
  wire _7645_;
  wire _7646_;
  wire _7647_;
  wire _7648_;
  wire _7649_;
  wire _7650_;
  wire _7651_;
  wire _7652_;
  wire _7653_;
  wire _7654_;
  wire _7655_;
  wire _7656_;
  wire _7657_;
  wire _7658_;
  wire _7659_;
  wire _7660_;
  wire _7661_;
  wire _7662_;
  wire _7663_;
  wire _7664_;
  wire _7665_;
  wire _7666_;
  wire _7667_;
  wire _7668_;
  wire _7669_;
  wire _7670_;
  wire _7671_;
  wire _7672_;
  wire _7673_;
  wire _7674_;
  wire _7675_;
  wire _7676_;
  wire _7677_;
  wire _7678_;
  wire _7679_;
  wire _7680_;
  wire _7681_;
  wire _7682_;
  wire _7683_;
  wire _7684_;
  wire _7685_;
  wire _7686_;
  wire _7687_;
  wire _7688_;
  wire _7689_;
  wire _7690_;
  wire _7691_;
  wire _7692_;
  wire _7693_;
  wire _7694_;
  wire _7695_;
  wire _7696_;
  wire _7697_;
  wire _7698_;
  wire _7699_;
  wire _7700_;
  wire _7701_;
  wire _7702_;
  wire _7703_;
  wire _7704_;
  wire _7705_;
  wire _7706_;
  wire _7707_;
  wire _7708_;
  wire _7709_;
  wire _7710_;
  wire _7711_;
  wire _7712_;
  wire _7713_;
  wire _7714_;
  wire _7715_;
  wire _7716_;
  wire _7717_;
  wire _7718_;
  wire _7719_;
  wire _7720_;
  wire _7721_;
  wire _7722_;
  wire _7723_;
  wire _7724_;
  wire _7725_;
  wire _7726_;
  wire _7727_;
  wire _7728_;
  wire _7729_;
  wire _7730_;
  wire _7731_;
  wire _7732_;
  wire _7733_;
  wire _7734_;
  wire _7735_;
  wire _7736_;
  wire _7737_;
  wire _7738_;
  wire _7739_;
  wire _7740_;
  wire _7741_;
  wire _7742_;
  wire _7743_;
  wire _7744_;
  wire _7745_;
  wire _7746_;
  wire _7747_;
  wire _7748_;
  wire _7749_;
  wire _7750_;
  wire _7751_;
  wire _7752_;
  wire _7753_;
  wire _7754_;
  wire _7755_;
  wire _7756_;
  wire _7757_;
  wire _7758_;
  wire _7759_;
  wire _7760_;
  wire _7761_;
  wire _7762_;
  wire _7763_;
  wire _7764_;
  wire _7765_;
  wire _7766_;
  wire _7767_;
  wire _7768_;
  wire _7769_;
  wire _7770_;
  wire _7771_;
  wire _7772_;
  wire _7773_;
  wire _7774_;
  wire _7775_;
  wire _7776_;
  wire _7777_;
  wire _7778_;
  wire _7779_;
  wire _7780_;
  wire _7781_;
  wire _7782_;
  wire _7783_;
  wire _7784_;
  wire _7785_;
  wire _7786_;
  wire _7787_;
  wire _7788_;
  wire _7789_;
  wire _7790_;
  wire _7791_;
  wire _7792_;
  wire _7793_;
  wire _7794_;
  wire _7795_;
  wire _7796_;
  wire _7797_;
  wire _7798_;
  wire _7799_;
  wire _7800_;
  wire _7801_;
  wire _7802_;
  wire _7803_;
  wire _7804_;
  wire _7805_;
  wire _7806_;
  wire _7807_;
  wire _7808_;
  wire _7809_;
  wire _7810_;
  wire _7811_;
  wire _7812_;
  wire _7813_;
  wire _7814_;
  wire _7815_;
  wire _7816_;
  wire _7817_;
  wire _7818_;
  wire _7819_;
  wire _7820_;
  wire _7821_;
  wire _7822_;
  wire _7823_;
  wire _7824_;
  wire _7825_;
  wire _7826_;
  wire _7827_;
  wire _7828_;
  wire _7829_;
  wire _7830_;
  wire _7831_;
  wire _7832_;
  wire _7833_;
  wire _7834_;
  wire _7835_;
  wire _7836_;
  wire _7837_;
  wire _7838_;
  wire _7839_;
  wire _7840_;
  wire _7841_;
  wire _7842_;
  wire _7843_;
  wire _7844_;
  wire _7845_;
  wire _7846_;
  wire _7847_;
  wire _7848_;
  wire _7849_;
  wire _7850_;
  wire _7851_;
  wire _7852_;
  wire _7853_;
  wire _7854_;
  wire _7855_;
  wire _7856_;
  wire _7857_;
  wire _7858_;
  wire _7859_;
  wire _7860_;
  wire _7861_;
  wire _7862_;
  wire _7863_;
  wire _7864_;
  wire _7865_;
  wire _7866_;
  wire _7867_;
  wire _7868_;
  wire _7869_;
  wire _7870_;
  wire _7871_;
  wire _7872_;
  wire _7873_;
  wire _7874_;
  wire _7875_;
  wire _7876_;
  wire _7877_;
  wire _7878_;
  wire _7879_;
  wire _7880_;
  wire _7881_;
  wire _7882_;
  wire _7883_;
  wire _7884_;
  wire _7885_;
  wire _7886_;
  wire _7887_;
  wire _7888_;
  wire _7889_;
  wire _7890_;
  wire _7891_;
  wire _7892_;
  wire _7893_;
  wire _7894_;
  wire _7895_;
  wire _7896_;
  wire _7897_;
  wire _7898_;
  wire _7899_;
  wire _7900_;
  wire _7901_;
  wire _7902_;
  wire _7903_;
  wire _7904_;
  wire _7905_;
  wire _7906_;
  wire _7907_;
  wire _7908_;
  wire _7909_;
  wire _7910_;
  wire _7911_;
  wire _7912_;
  wire _7913_;
  wire _7914_;
  wire _7915_;
  wire _7916_;
  wire _7917_;
  wire _7918_;
  wire _7919_;
  wire _7920_;
  wire _7921_;
  wire _7922_;
  wire _7923_;
  wire _7924_;
  wire _7925_;
  wire _7926_;
  wire _7927_;
  wire _7928_;
  wire _7929_;
  wire _7930_;
  wire _7931_;
  wire _7932_;
  wire _7933_;
  wire _7934_;
  wire _7935_;
  wire _7936_;
  wire _7937_;
  wire _7938_;
  wire _7939_;
  wire _7940_;
  wire _7941_;
  wire _7942_;
  wire _7943_;
  wire _7944_;
  wire _7945_;
  wire _7946_;
  wire _7947_;
  wire _7948_;
  wire _7949_;
  wire _7950_;
  wire _7951_;
  wire _7952_;
  wire _7953_;
  wire _7954_;
  wire _7955_;
  wire _7956_;
  wire _7957_;
  wire _7958_;
  wire _7959_;
  wire _7960_;
  wire _7961_;
  wire _7962_;
  wire _7963_;
  wire _7964_;
  wire _7965_;
  wire _7966_;
  wire _7967_;
  wire _7968_;
  wire _7969_;
  wire _7970_;
  wire _7971_;
  wire _7972_;
  wire _7973_;
  wire _7974_;
  wire _7975_;
  wire _7976_;
  wire _7977_;
  wire _7978_;
  wire _7979_;
  wire _7980_;
  wire _7981_;
  wire _7982_;
  wire _7983_;
  wire _7984_;
  wire _7985_;
  wire _7986_;
  wire _7987_;
  wire _7988_;
  wire _7989_;
  wire _7990_;
  wire _7991_;
  wire _7992_;
  wire _7993_;
  wire _7994_;
  wire _7995_;
  wire _7996_;
  wire _7997_;
  wire _7998_;
  wire _7999_;
  wire _8000_;
  wire _8001_;
  wire _8002_;
  wire _8003_;
  wire _8004_;
  wire _8005_;
  wire _8006_;
  wire _8007_;
  wire _8008_;
  wire _8009_;
  wire _8010_;
  wire _8011_;
  wire _8012_;
  wire _8013_;
  wire _8014_;
  wire _8015_;
  wire _8016_;
  wire _8017_;
  wire _8018_;
  wire _8019_;
  wire _8020_;
  wire _8021_;
  wire _8022_;
  wire _8023_;
  wire _8024_;
  wire _8025_;
  wire _8026_;
  wire _8027_;
  wire _8028_;
  wire _8029_;
  wire _8030_;
  wire _8031_;
  wire _8032_;
  wire _8033_;
  wire _8034_;
  wire _8035_;
  wire _8036_;
  wire _8037_;
  wire _8038_;
  wire _8039_;
  wire _8040_;
  wire _8041_;
  wire _8042_;
  wire _8043_;
  wire _8044_;
  wire _8045_;
  wire _8046_;
  wire _8047_;
  wire _8048_;
  wire _8049_;
  wire _8050_;
  wire _8051_;
  wire _8052_;
  wire _8053_;
  wire _8054_;
  wire _8055_;
  wire _8056_;
  wire _8057_;
  wire _8058_;
  wire _8059_;
  wire _8060_;
  wire _8061_;
  wire _8062_;
  wire _8063_;
  wire _8064_;
  wire _8065_;
  wire _8066_;
  wire _8067_;
  wire _8068_;
  wire _8069_;
  wire _8070_;
  wire _8071_;
  wire _8072_;
  wire _8073_;
  wire _8074_;
  wire _8075_;
  wire _8076_;
  wire _8077_;
  wire _8078_;
  wire _8079_;
  wire _8080_;
  wire _8081_;
  wire _8082_;
  wire _8083_;
  wire _8084_;
  wire _8085_;
  wire _8086_;
  wire _8087_;
  wire _8088_;
  wire _8089_;
  wire _8090_;
  wire _8091_;
  wire _8092_;
  wire _8093_;
  wire _8094_;
  wire _8095_;
  wire _8096_;
  wire _8097_;
  wire _8098_;
  wire _8099_;
  wire _8100_;
  wire _8101_;
  wire _8102_;
  wire _8103_;
  wire _8104_;
  wire _8105_;
  wire _8106_;
  wire _8107_;
  wire _8108_;
  wire _8109_;
  wire _8110_;
  wire _8111_;
  wire _8112_;
  wire _8113_;
  wire _8114_;
  wire _8115_;
  wire _8116_;
  wire _8117_;
  wire _8118_;
  wire _8119_;
  wire _8120_;
  wire _8121_;
  wire _8122_;
  wire _8123_;
  wire _8124_;
  wire _8125_;
  wire _8126_;
  wire _8127_;
  wire _8128_;
  wire _8129_;
  wire _8130_;
  wire _8131_;
  wire _8132_;
  wire _8133_;
  wire _8134_;
  wire _8135_;
  wire _8136_;
  wire _8137_;
  wire _8138_;
  wire _8139_;
  wire _8140_;
  wire _8141_;
  wire _8142_;
  wire _8143_;
  wire _8144_;
  wire _8145_;
  wire _8146_;
  wire _8147_;
  wire _8148_;
  wire _8149_;
  wire _8150_;
  wire _8151_;
  wire _8152_;
  wire _8153_;
  wire _8154_;
  wire _8155_;
  wire _8156_;
  wire _8157_;
  wire _8158_;
  wire _8159_;
  wire _8160_;
  wire _8161_;
  wire _8162_;
  wire _8163_;
  wire _8164_;
  wire _8165_;
  wire _8166_;
  wire _8167_;
  wire _8168_;
  wire _8169_;
  wire _8170_;
  wire _8171_;
  wire _8172_;
  wire _8173_;
  wire _8174_;
  wire _8175_;
  wire _8176_;
  wire _8177_;
  wire _8178_;
  wire _8179_;
  wire _8180_;
  wire _8181_;
  wire _8182_;
  wire _8183_;
  wire _8184_;
  wire _8185_;
  wire _8186_;
  wire _8187_;
  wire _8188_;
  wire _8189_;
  wire _8190_;
  wire _8191_;
  wire _8192_;
  wire _8193_;
  wire _8194_;
  wire _8195_;
  wire _8196_;
  wire _8197_;
  wire _8198_;
  wire _8199_;
  wire _8200_;
  wire _8201_;
  wire _8202_;
  wire _8203_;
  wire _8204_;
  wire _8205_;
  wire _8206_;
  wire _8207_;
  wire _8208_;
  wire _8209_;
  wire _8210_;
  wire _8211_;
  wire _8212_;
  wire _8213_;
  wire _8214_;
  wire _8215_;
  wire _8216_;
  wire _8217_;
  wire _8218_;
  wire _8219_;
  wire _8220_;
  wire _8221_;
  wire _8222_;
  wire _8223_;
  wire _8224_;
  wire _8225_;
  wire _8226_;
  wire _8227_;
  wire _8228_;
  wire _8229_;
  wire _8230_;
  wire _8231_;
  wire _8232_;
  wire _8233_;
  wire _8234_;
  wire _8235_;
  wire _8236_;
  wire _8237_;
  wire _8238_;
  wire _8239_;
  wire _8240_;
  wire _8241_;
  wire _8242_;
  wire _8243_;
  wire _8244_;
  wire _8245_;
  wire _8246_;
  wire _8247_;
  wire _8248_;
  wire _8249_;
  wire _8250_;
  wire _8251_;
  wire _8252_;
  wire _8253_;
  wire _8254_;
  wire _8255_;
  wire _8256_;
  wire _8257_;
  wire _8258_;
  wire _8259_;
  wire _8260_;
  wire _8261_;
  wire _8262_;
  wire _8263_;
  wire _8264_;
  wire _8265_;
  wire _8266_;
  wire _8267_;
  wire _8268_;
  wire _8269_;
  wire _8270_;
  wire _8271_;
  wire _8272_;
  wire _8273_;
  wire _8274_;
  wire _8275_;
  wire _8276_;
  wire _8277_;
  wire _8278_;
  wire _8279_;
  wire _8280_;
  wire _8281_;
  wire _8282_;
  wire _8283_;
  wire _8284_;
  wire _8285_;
  wire _8286_;
  wire _8287_;
  wire _8288_;
  wire _8289_;
  wire _8290_;
  wire _8291_;
  wire _8292_;
  wire _8293_;
  wire _8294_;
  wire _8295_;
  wire _8296_;
  wire _8297_;
  wire _8298_;
  wire _8299_;
  wire _8300_;
  wire _8301_;
  wire _8302_;
  wire _8303_;
  wire _8304_;
  wire _8305_;
  wire _8306_;
  wire _8307_;
  wire _8308_;
  wire _8309_;
  wire _8310_;
  wire _8311_;
  wire _8312_;
  wire _8313_;
  wire _8314_;
  wire _8315_;
  wire _8316_;
  wire _8317_;
  wire _8318_;
  wire _8319_;
  wire _8320_;
  wire _8321_;
  wire _8322_;
  wire _8323_;
  wire _8324_;
  wire _8325_;
  wire _8326_;
  wire _8327_;
  wire _8328_;
  wire _8329_;
  wire _8330_;
  wire _8331_;
  wire _8332_;
  wire _8333_;
  wire _8334_;
  wire _8335_;
  wire _8336_;
  wire _8337_;
  wire _8338_;
  wire _8339_;
  wire _8340_;
  wire _8341_;
  wire _8342_;
  wire _8343_;
  wire _8344_;
  wire _8345_;
  wire _8346_;
  wire _8347_;
  wire _8348_;
  wire _8349_;
  wire _8350_;
  wire _8351_;
  wire _8352_;
  wire _8353_;
  wire _8354_;
  wire _8355_;
  wire _8356_;
  wire _8357_;
  wire _8358_;
  wire _8359_;
  wire _8360_;
  wire _8361_;
  wire _8362_;
  wire _8363_;
  wire _8364_;
  wire _8365_;
  wire _8366_;
  wire _8367_;
  wire _8368_;
  wire _8369_;
  wire _8370_;
  wire _8371_;
  wire _8372_;
  wire _8373_;
  wire _8374_;
  wire _8375_;
  wire _8376_;
  wire _8377_;
  wire _8378_;
  wire _8379_;
  wire _8380_;
  wire _8381_;
  wire _8382_;
  wire _8383_;
  wire _8384_;
  wire _8385_;
  wire _8386_;
  wire _8387_;
  wire _8388_;
  wire _8389_;
  wire _8390_;
  wire _8391_;
  wire _8392_;
  wire _8393_;
  wire _8394_;
  wire _8395_;
  wire _8396_;
  wire _8397_;
  wire _8398_;
  wire _8399_;
  wire _8400_;
  wire _8401_;
  wire _8402_;
  wire _8403_;
  wire _8404_;
  wire _8405_;
  wire _8406_;
  wire _8407_;
  wire _8408_;
  wire _8409_;
  wire _8410_;
  wire _8411_;
  wire _8412_;
  wire _8413_;
  wire _8414_;
  wire _8415_;
  wire _8416_;
  wire _8417_;
  wire _8418_;
  wire _8419_;
  wire _8420_;
  wire _8421_;
  wire _8422_;
  wire _8423_;
  wire _8424_;
  wire _8425_;
  wire _8426_;
  wire _8427_;
  wire _8428_;
  wire _8429_;
  wire _8430_;
  wire _8431_;
  wire _8432_;
  wire _8433_;
  wire _8434_;
  wire _8435_;
  wire _8436_;
  wire _8437_;
  wire _8438_;
  wire _8439_;
  wire _8440_;
  wire _8441_;
  wire _8442_;
  wire _8443_;
  wire _8444_;
  wire _8445_;
  wire _8446_;
  wire _8447_;
  wire _8448_;
  wire _8449_;
  wire _8450_;
  wire _8451_;
  wire _8452_;
  wire _8453_;
  wire _8454_;
  wire _8455_;
  wire _8456_;
  wire _8457_;
  wire _8458_;
  wire _8459_;
  wire _8460_;
  wire _8461_;
  wire _8462_;
  wire _8463_;
  wire _8464_;
  wire _8465_;
  wire _8466_;
  wire _8467_;
  wire _8468_;
  wire _8469_;
  wire _8470_;
  wire _8471_;
  wire _8472_;
  wire _8473_;
  wire _8474_;
  wire _8475_;
  wire _8476_;
  wire _8477_;
  wire _8478_;
  wire _8479_;
  wire _8480_;
  wire _8481_;
  wire _8482_;
  wire _8483_;
  wire _8484_;
  wire _8485_;
  wire _8486_;
  wire _8487_;
  wire _8488_;
  wire _8489_;
  wire _8490_;
  wire _8491_;
  wire _8492_;
  wire _8493_;
  wire _8494_;
  wire _8495_;
  wire _8496_;
  wire _8497_;
  wire _8498_;
  wire _8499_;
  wire _8500_;
  wire _8501_;
  wire _8502_;
  wire _8503_;
  wire _8504_;
  wire _8505_;
  wire _8506_;
  wire _8507_;
  wire _8508_;
  wire _8509_;
  wire _8510_;
  wire _8511_;
  wire _8512_;
  wire _8513_;
  wire _8514_;
  wire _8515_;
  wire _8516_;
  wire _8517_;
  wire _8518_;
  wire _8519_;
  wire _8520_;
  wire _8521_;
  wire _8522_;
  wire _8523_;
  wire _8524_;
  wire _8525_;
  wire _8526_;
  wire _8527_;
  wire _8528_;
  wire _8529_;
  wire _8530_;
  wire _8531_;
  wire _8532_;
  wire _8533_;
  wire _8534_;
  wire _8535_;
  wire _8536_;
  wire _8537_;
  wire _8538_;
  wire _8539_;
  wire _8540_;
  wire _8541_;
  wire _8542_;
  wire _8543_;
  wire _8544_;
  wire _8545_;
  wire _8546_;
  wire _8547_;
  wire _8548_;
  wire _8549_;
  wire _8550_;
  wire _8551_;
  wire _8552_;
  wire _8553_;
  wire _8554_;
  wire _8555_;
  wire _8556_;
  wire _8557_;
  wire _8558_;
  wire _8559_;
  wire _8560_;
  wire _8561_;
  wire _8562_;
  wire _8563_;
  wire _8564_;
  wire _8565_;
  wire _8566_;
  wire _8567_;
  wire _8568_;
  wire _8569_;
  wire _8570_;
  wire _8571_;
  wire _8572_;
  wire _8573_;
  wire _8574_;
  wire _8575_;
  wire _8576_;
  wire _8577_;
  wire _8578_;
  wire _8579_;
  wire _8580_;
  wire _8581_;
  wire _8582_;
  wire _8583_;
  wire _8584_;
  wire _8585_;
  wire _8586_;
  wire _8587_;
  wire _8588_;
  wire _8589_;
  wire _8590_;
  wire _8591_;
  wire _8592_;
  wire _8593_;
  wire _8594_;
  wire _8595_;
  wire _8596_;
  wire _8597_;
  wire _8598_;
  wire _8599_;
  wire _8600_;
  wire _8601_;
  wire _8602_;
  wire _8603_;
  wire _8604_;
  wire _8605_;
  wire _8606_;
  wire _8607_;
  wire _8608_;
  wire _8609_;
  wire _8610_;
  wire _8611_;
  wire _8612_;
  wire _8613_;
  wire _8614_;
  wire _8615_;
  wire _8616_;
  wire _8617_;
  wire _8618_;
  wire _8619_;
  wire _8620_;
  wire _8621_;
  wire _8622_;
  wire _8623_;
  wire _8624_;
  wire _8625_;
  wire _8626_;
  wire _8627_;
  wire _8628_;
  wire _8629_;
  wire _8630_;
  wire _8631_;
  wire _8632_;
  wire _8633_;
  wire _8634_;
  wire _8635_;
  wire _8636_;
  wire _8637_;
  wire _8638_;
  wire _8639_;
  wire _8640_;
  wire _8641_;
  wire _8642_;
  wire _8643_;
  wire _8644_;
  wire _8645_;
  wire _8646_;
  wire _8647_;
  wire _8648_;
  wire _8649_;
  wire _8650_;
  wire _8651_;
  wire _8652_;
  wire _8653_;
  wire _8654_;
  wire _8655_;
  wire _8656_;
  wire _8657_;
  wire _8658_;
  wire _8659_;
  wire _8660_;
  wire _8661_;
  wire _8662_;
  wire _8663_;
  wire _8664_;
  wire _8665_;
  wire _8666_;
  wire _8667_;
  wire _8668_;
  wire _8669_;
  wire _8670_;
  wire _8671_;
  wire _8672_;
  wire _8673_;
  wire _8674_;
  wire _8675_;
  wire _8676_;
  wire _8677_;
  wire _8678_;
  wire _8679_;
  wire _8680_;
  wire _8681_;
  wire _8682_;
  wire _8683_;
  wire _8684_;
  wire _8685_;
  wire _8686_;
  wire _8687_;
  wire _8688_;
  wire _8689_;
  wire _8690_;
  wire _8691_;
  wire _8692_;
  wire _8693_;
  wire _8694_;
  wire _8695_;
  wire _8696_;
  wire _8697_;
  wire _8698_;
  wire _8699_;
  wire _8700_;
  wire _8701_;
  wire _8702_;
  wire _8703_;
  wire _8704_;
  wire _8705_;
  wire _8706_;
  wire _8707_;
  wire _8708_;
  wire _8709_;
  wire _8710_;
  wire _8711_;
  wire _8712_;
  wire _8713_;
  wire _8714_;
  wire _8715_;
  wire _8716_;
  wire _8717_;
  wire _8718_;
  wire _8719_;
  wire _8720_;
  wire _8721_;
  wire _8722_;
  wire _8723_;
  wire _8724_;
  wire _8725_;
  wire _8726_;
  wire _8727_;
  wire _8728_;
  wire _8729_;
  wire _8730_;
  wire _8731_;
  wire _8732_;
  wire _8733_;
  wire _8734_;
  wire _8735_;
  wire _8736_;
  wire _8737_;
  wire _8738_;
  wire _8739_;
  wire _8740_;
  wire _8741_;
  wire _8742_;
  wire _8743_;
  wire _8744_;
  wire _8745_;
  wire _8746_;
  wire _8747_;
  wire _8748_;
  wire _8749_;
  wire _8750_;
  wire _8751_;
  wire _8752_;
  wire _8753_;
  wire _8754_;
  wire _8755_;
  wire _8756_;
  wire _8757_;
  wire _8758_;
  wire _8759_;
  wire _8760_;
  wire _8761_;
  wire _8762_;
  wire _8763_;
  wire _8764_;
  wire _8765_;
  wire _8766_;
  wire _8767_;
  wire _8768_;
  wire _8769_;
  wire _8770_;
  wire _8771_;
  wire _8772_;
  wire _8773_;
  wire _8774_;
  wire _8775_;
  wire _8776_;
  wire _8777_;
  wire _8778_;
  wire _8779_;
  wire _8780_;
  wire _8781_;
  wire _8782_;
  wire _8783_;
  wire _8784_;
  wire _8785_;
  wire _8786_;
  wire _8787_;
  wire _8788_;
  wire _8789_;
  wire _8790_;
  wire _8791_;
  wire _8792_;
  wire _8793_;
  wire _8794_;
  wire _8795_;
  wire _8796_;
  wire _8797_;
  wire _8798_;
  wire _8799_;
  wire _8800_;
  wire _8801_;
  wire _8802_;
  wire _8803_;
  wire _8804_;
  wire _8805_;
  wire _8806_;
  wire _8807_;
  wire _8808_;
  wire _8809_;
  wire _8810_;
  wire _8811_;
  wire _8812_;
  wire _8813_;
  wire _8814_;
  wire _8815_;
  wire _8816_;
  wire _8817_;
  wire _8818_;
  wire _8819_;
  wire _8820_;
  wire _8821_;
  wire _8822_;
  wire _8823_;
  wire _8824_;
  wire _8825_;
  wire _8826_;
  wire _8827_;
  wire _8828_;
  wire _8829_;
  wire _8830_;
  wire _8831_;
  wire _8832_;
  wire _8833_;
  wire _8834_;
  wire _8835_;
  wire _8836_;
  wire _8837_;
  wire _8838_;
  wire _8839_;
  wire _8840_;
  wire _8841_;
  wire _8842_;
  wire _8843_;
  wire _8844_;
  wire _8845_;
  wire _8846_;
  wire _8847_;
  wire _8848_;
  wire _8849_;
  wire _8850_;
  wire _8851_;
  wire _8852_;
  wire _8853_;
  wire _8854_;
  wire _8855_;
  wire _8856_;
  wire _8857_;
  wire _8858_;
  wire _8859_;
  wire _8860_;
  wire _8861_;
  wire _8862_;
  wire _8863_;
  wire _8864_;
  wire _8865_;
  wire _8866_;
  wire _8867_;
  wire _8868_;
  wire _8869_;
  wire _8870_;
  wire _8871_;
  wire _8872_;
  wire _8873_;
  wire _8874_;
  wire _8875_;
  wire _8876_;
  wire _8877_;
  wire _8878_;
  wire _8879_;
  wire _8880_;
  wire _8881_;
  wire _8882_;
  wire _8883_;
  wire _8884_;
  wire _8885_;
  wire _8886_;
  wire _8887_;
  wire _8888_;
  wire _8889_;
  wire _8890_;
  wire _8891_;
  wire _8892_;
  wire _8893_;
  wire _8894_;
  wire _8895_;
  wire _8896_;
  wire _8897_;
  wire _8898_;
  wire _8899_;
  wire _8900_;
  wire _8901_;
  wire _8902_;
  wire _8903_;
  wire _8904_;
  wire _8905_;
  wire _8906_;
  wire _8907_;
  wire _8908_;
  wire _8909_;
  wire _8910_;
  wire _8911_;
  wire _8912_;
  wire _8913_;
  wire _8914_;
  wire _8915_;
  wire _8916_;
  wire _8917_;
  wire _8918_;
  wire _8919_;
  wire _8920_;
  wire _8921_;
  wire _8922_;
  wire _8923_;
  wire _8924_;
  wire _8925_;
  wire _8926_;
  wire _8927_;
  wire _8928_;
  wire _8929_;
  wire _8930_;
  wire _8931_;
  wire _8932_;
  wire _8933_;
  wire _8934_;
  wire _8935_;
  wire _8936_;
  wire _8937_;
  wire _8938_;
  wire _8939_;
  wire _8940_;
  wire _8941_;
  wire _8942_;
  wire _8943_;
  wire _8944_;
  wire _8945_;
  wire _8946_;
  wire _8947_;
  wire _8948_;
  wire _8949_;
  wire _8950_;
  wire _8951_;
  wire _8952_;
  wire _8953_;
  wire _8954_;
  wire _8955_;
  wire _8956_;
  wire _8957_;
  wire _8958_;
  wire _8959_;
  wire _8960_;
  wire _8961_;
  wire _8962_;
  wire _8963_;
  wire _8964_;
  wire _8965_;
  wire _8966_;
  wire _8967_;
  wire _8968_;
  wire _8969_;
  wire _8970_;
  wire _8971_;
  wire _8972_;
  wire _8973_;
  wire _8974_;
  wire _8975_;
  wire _8976_;
  wire _8977_;
  wire _8978_;
  wire _8979_;
  wire _8980_;
  wire _8981_;
  wire _8982_;
  wire _8983_;
  wire _8984_;
  wire _8985_;
  wire _8986_;
  wire _8987_;
  wire _8988_;
  wire _8989_;
  wire _8990_;
  wire _8991_;
  wire _8992_;
  wire _8993_;
  wire _8994_;
  wire _8995_;
  wire _8996_;
  wire _8997_;
  wire _8998_;
  wire _8999_;
  wire _9000_;
  wire _9001_;
  wire _9002_;
  wire _9003_;
  wire _9004_;
  wire _9005_;
  wire _9006_;
  wire _9007_;
  wire _9008_;
  wire _9009_;
  wire _9010_;
  wire _9011_;
  wire _9012_;
  wire _9013_;
  wire _9014_;
  wire _9015_;
  wire _9016_;
  wire _9017_;
  wire _9018_;
  wire _9019_;
  wire _9020_;
  wire _9021_;
  wire _9022_;
  wire _9023_;
  wire _9024_;
  wire _9025_;
  wire _9026_;
  wire _9027_;
  wire _9028_;
  wire _9029_;
  wire _9030_;
  wire _9031_;
  wire _9032_;
  wire _9033_;
  wire _9034_;
  wire _9035_;
  wire _9036_;
  wire _9037_;
  wire _9038_;
  wire _9039_;
  wire _9040_;
  wire _9041_;
  wire _9042_;
  wire _9043_;
  wire _9044_;
  wire _9045_;
  wire _9046_;
  wire _9047_;
  wire _9048_;
  wire _9049_;
  wire _9050_;
  wire _9051_;
  wire _9052_;
  wire _9053_;
  wire _9054_;
  wire _9055_;
  wire _9056_;
  wire _9057_;
  wire _9058_;
  wire _9059_;
  wire _9060_;
  wire _9061_;
  wire _9062_;
  wire _9063_;
  wire _9064_;
  wire _9065_;
  wire _9066_;
  wire _9067_;
  wire _9068_;
  wire _9069_;
  wire _9070_;
  wire _9071_;
  wire _9072_;
  wire _9073_;
  wire _9074_;
  wire _9075_;
  wire _9076_;
  wire _9077_;
  wire _9078_;
  wire _9079_;
  wire _9080_;
  wire _9081_;
  wire _9082_;
  wire _9083_;
  wire _9084_;
  wire _9085_;
  wire _9086_;
  wire _9087_;
  wire _9088_;
  wire _9089_;
  wire _9090_;
  wire _9091_;
  wire _9092_;
  wire _9093_;
  wire _9094_;
  wire _9095_;
  wire _9096_;
  wire _9097_;
  wire _9098_;
  wire _9099_;
  wire _9100_;
  wire _9101_;
  wire _9102_;
  wire _9103_;
  wire _9104_;
  wire _9105_;
  wire _9106_;
  wire _9107_;
  wire _9108_;
  wire _9109_;
  wire _9110_;
  wire _9111_;
  wire _9112_;
  wire _9113_;
  wire _9114_;
  wire _9115_;
  wire _9116_;
  wire _9117_;
  wire _9118_;
  wire _9119_;
  wire _9120_;
  wire _9121_;
  wire _9122_;
  wire _9123_;
  wire _9124_;
  wire _9125_;
  wire _9126_;
  wire _9127_;
  wire _9128_;
  wire _9129_;
  wire _9130_;
  wire _9131_;
  wire _9132_;
  wire _9133_;
  wire _9134_;
  wire _9135_;
  wire _9136_;
  wire _9137_;
  wire _9138_;
  wire _9139_;
  wire _9140_;
  wire _9141_;
  wire _9142_;
  wire _9143_;
  wire _9144_;
  wire _9145_;
  wire _9146_;
  wire _9147_;
  wire _9148_;
  wire _9149_;
  wire _9150_;
  wire _9151_;
  wire _9152_;
  wire _9153_;
  wire _9154_;
  wire _9155_;
  wire _9156_;
  wire _9157_;
  wire _9158_;
  wire _9159_;
  wire _9160_;
  wire _9161_;
  wire _9162_;
  wire _9163_;
  wire _9164_;
  wire _9165_;
  wire _9166_;
  wire _9167_;
  wire _9168_;
  wire _9169_;
  wire _9170_;
  wire _9171_;
  wire _9172_;
  wire _9173_;
  wire _9174_;
  wire _9175_;
  wire _9176_;
  wire _9177_;
  wire _9178_;
  wire _9179_;
  wire _9180_;
  wire _9181_;
  wire _9182_;
  wire _9183_;
  wire _9184_;
  wire _9185_;
  wire _9186_;
  wire _9187_;
  wire _9188_;
  wire _9189_;
  wire _9190_;
  wire _9191_;
  wire _9192_;
  wire _9193_;
  wire _9194_;
  wire _9195_;
  wire _9196_;
  wire _9197_;
  wire _9198_;
  wire _9199_;
  wire _9200_;
  wire _9201_;
  wire _9202_;
  wire _9203_;
  wire _9204_;
  wire _9205_;
  wire _9206_;
  wire _9207_;
  wire _9208_;
  wire _9209_;
  wire _9210_;
  wire _9211_;
  wire _9212_;
  wire _9213_;
  wire _9214_;
  wire _9215_;
  wire _9216_;
  wire _9217_;
  wire _9218_;
  wire _9219_;
  wire _9220_;
  wire _9221_;
  wire _9222_;
  wire _9223_;
  wire _9224_;
  wire _9225_;
  wire _9226_;
  wire _9227_;
  wire _9228_;
  wire _9229_;
  wire _9230_;
  wire _9231_;
  wire _9232_;
  wire _9233_;
  wire _9234_;
  wire _9235_;
  wire _9236_;
  wire _9237_;
  wire _9238_;
  wire _9239_;
  wire _9240_;
  wire _9241_;
  wire _9242_;
  wire _9243_;
  wire _9244_;
  wire _9245_;
  wire _9246_;
  wire _9247_;
  wire _9248_;
  wire _9249_;
  wire _9250_;
  wire _9251_;
  wire _9252_;
  wire _9253_;
  wire _9254_;
  wire _9255_;
  wire _9256_;
  wire _9257_;
  wire _9258_;
  wire _9259_;
  wire _9260_;
  wire _9261_;
  wire _9262_;
  wire _9263_;
  wire _9264_;
  wire _9265_;
  wire _9266_;
  wire _9267_;
  wire _9268_;
  wire _9269_;
  wire _9270_;
  wire _9271_;
  wire _9272_;
  wire _9273_;
  wire _9274_;
  wire _9275_;
  wire _9276_;
  wire _9277_;
  wire _9278_;
  wire _9279_;
  wire _9280_;
  wire _9281_;
  wire _9282_;
  wire _9283_;
  wire _9284_;
  wire _9285_;
  wire _9286_;
  wire _9287_;
  wire _9288_;
  wire _9289_;
  wire _9290_;
  wire _9291_;
  wire _9292_;
  wire _9293_;
  wire _9294_;
  wire _9295_;
  wire _9296_;
  wire _9297_;
  wire alu_valid_id_ex;
  wire alu_valid_id_ex_t0;
  wire alu_valid_id_ex_t1;
  wire [3:0] \amo_req.amo_op ;
  wire [63:0] \amo_req.operand_a ;
  wire [63:0] \amo_req.operand_b ;
  wire \amo_req.req ;
  wire [1:0] \amo_req.size ;
  wire \amo_resp.ack ;
  wire \amo_resp.ack_t0 ;
  wire \amo_resp.ack_t1 ;
  wire [63:0] \amo_resp.result ;
  wire [63:0] \amo_resp.result_t0 ;
  wire [63:0] \amo_resp.result_t1 ;
  wire amo_valid_commit;
  wire amo_valid_commit_t0;
  wire amo_valid_commit_t1;
  wire [15:0] asid_csr_ex;
  wire [15:0] asid_csr_ex_t0;
  wire [15:0] asid_csr_ex_t1;
  wire [63:0] boot_addr_i;
  wire [63:0] boot_addr_i_t0;
  wire [63:0] boot_addr_i_t1;
  wire [2:0] \branch_predict_id_ex.cf ;
  wire [2:0] \branch_predict_id_ex.cf_t0 ;
  wire [2:0] \branch_predict_id_ex.cf_t1 ;
  wire [63:0] \branch_predict_id_ex.predict_address ;
  wire [63:0] \branch_predict_id_ex.predict_address_t0 ;
  wire [63:0] \branch_predict_id_ex.predict_address_t1 ;
  wire branch_valid_id_ex;
  wire branch_valid_id_ex_t0;
  wire branch_valid_id_ex_t1;
  wire [1:0] commit_ack;
  wire [1:0] commit_ack_t0;
  wire [1:0] commit_ack_t1;
  wire [2:0] \commit_instr_id_commit[0].bp.cf ;
  wire [2:0] \commit_instr_id_commit[0].bp.cf_t0 ;
  wire [2:0] \commit_instr_id_commit[0].bp.cf_t1 ;
  wire [63:0] \commit_instr_id_commit[0].bp.predict_address ;
  wire [63:0] \commit_instr_id_commit[0].bp.predict_address_t0 ;
  wire [63:0] \commit_instr_id_commit[0].bp.predict_address_t1 ;
  wire [63:0] \commit_instr_id_commit[0].ex.cause ;
  wire [63:0] \commit_instr_id_commit[0].ex.cause_t0 ;
  wire [63:0] \commit_instr_id_commit[0].ex.cause_t1 ;
  wire [63:0] \commit_instr_id_commit[0].ex.tval ;
  wire [63:0] \commit_instr_id_commit[0].ex.tval_t0 ;
  wire [63:0] \commit_instr_id_commit[0].ex.tval_t1 ;
  wire \commit_instr_id_commit[0].ex.valid ;
  wire \commit_instr_id_commit[0].ex.valid_t0 ;
  wire \commit_instr_id_commit[0].ex.valid_t1 ;
  wire [3:0] \commit_instr_id_commit[0].fu ;
  wire [3:0] \commit_instr_id_commit[0].fu_t0 ;
  wire [3:0] \commit_instr_id_commit[0].fu_t1 ;
  wire \commit_instr_id_commit[0].is_compressed ;
  wire \commit_instr_id_commit[0].is_compressed_t0 ;
  wire \commit_instr_id_commit[0].is_compressed_t1 ;
  wire [6:0] \commit_instr_id_commit[0].op ;
  wire [6:0] \commit_instr_id_commit[0].op_t0 ;
  wire [6:0] \commit_instr_id_commit[0].op_t1 ;
  wire [63:0] \commit_instr_id_commit[0].pc ;
  wire [63:0] \commit_instr_id_commit[0].pc_t0 ;
  wire [63:0] \commit_instr_id_commit[0].pc_t1 ;
  wire [5:0] \commit_instr_id_commit[0].rd ;
  wire [5:0] \commit_instr_id_commit[0].rd_t0 ;
  wire [5:0] \commit_instr_id_commit[0].rd_t1 ;
  wire [63:0] \commit_instr_id_commit[0].result ;
  wire [63:0] \commit_instr_id_commit[0].result_t0 ;
  wire [63:0] \commit_instr_id_commit[0].result_t1 ;
  wire [5:0] \commit_instr_id_commit[0].rs1 ;
  wire [5:0] \commit_instr_id_commit[0].rs1_t0 ;
  wire [5:0] \commit_instr_id_commit[0].rs1_t1 ;
  wire [5:0] \commit_instr_id_commit[0].rs2 ;
  wire [5:0] \commit_instr_id_commit[0].rs2_t0 ;
  wire [5:0] \commit_instr_id_commit[0].rs2_t1 ;
  wire [1:0] \commit_instr_id_commit[0].trans_id ;
  wire [1:0] \commit_instr_id_commit[0].trans_id_t0 ;
  wire [1:0] \commit_instr_id_commit[0].trans_id_t1 ;
  wire \commit_instr_id_commit[0].use_imm ;
  wire \commit_instr_id_commit[0].use_imm_t0 ;
  wire \commit_instr_id_commit[0].use_imm_t1 ;
  wire \commit_instr_id_commit[0].use_pc ;
  wire \commit_instr_id_commit[0].use_pc_t0 ;
  wire \commit_instr_id_commit[0].use_pc_t1 ;
  wire \commit_instr_id_commit[0].use_zimm ;
  wire \commit_instr_id_commit[0].use_zimm_t0 ;
  wire \commit_instr_id_commit[0].use_zimm_t1 ;
  wire \commit_instr_id_commit[0].valid ;
  wire \commit_instr_id_commit[0].valid_t0 ;
  wire \commit_instr_id_commit[0].valid_t1 ;
  wire [2:0] \commit_instr_id_commit[1].bp.cf ;
  wire [2:0] \commit_instr_id_commit[1].bp.cf_t0 ;
  wire [2:0] \commit_instr_id_commit[1].bp.cf_t1 ;
  wire [63:0] \commit_instr_id_commit[1].bp.predict_address ;
  wire [63:0] \commit_instr_id_commit[1].bp.predict_address_t0 ;
  wire [63:0] \commit_instr_id_commit[1].bp.predict_address_t1 ;
  wire [63:0] \commit_instr_id_commit[1].ex.cause ;
  wire [63:0] \commit_instr_id_commit[1].ex.cause_t0 ;
  wire [63:0] \commit_instr_id_commit[1].ex.cause_t1 ;
  wire [63:0] \commit_instr_id_commit[1].ex.tval ;
  wire [63:0] \commit_instr_id_commit[1].ex.tval_t0 ;
  wire [63:0] \commit_instr_id_commit[1].ex.tval_t1 ;
  wire \commit_instr_id_commit[1].ex.valid ;
  wire \commit_instr_id_commit[1].ex.valid_t0 ;
  wire \commit_instr_id_commit[1].ex.valid_t1 ;
  wire [3:0] \commit_instr_id_commit[1].fu ;
  wire [3:0] \commit_instr_id_commit[1].fu_t0 ;
  wire [3:0] \commit_instr_id_commit[1].fu_t1 ;
  wire \commit_instr_id_commit[1].is_compressed ;
  wire \commit_instr_id_commit[1].is_compressed_t0 ;
  wire \commit_instr_id_commit[1].is_compressed_t1 ;
  wire [6:0] \commit_instr_id_commit[1].op ;
  wire [6:0] \commit_instr_id_commit[1].op_t0 ;
  wire [6:0] \commit_instr_id_commit[1].op_t1 ;
  wire [63:0] \commit_instr_id_commit[1].pc ;
  wire [63:0] \commit_instr_id_commit[1].pc_t0 ;
  wire [63:0] \commit_instr_id_commit[1].pc_t1 ;
  wire [5:0] \commit_instr_id_commit[1].rd ;
  wire [5:0] \commit_instr_id_commit[1].rd_t0 ;
  wire [5:0] \commit_instr_id_commit[1].rd_t1 ;
  wire [63:0] \commit_instr_id_commit[1].result ;
  wire [63:0] \commit_instr_id_commit[1].result_t0 ;
  wire [63:0] \commit_instr_id_commit[1].result_t1 ;
  wire [5:0] \commit_instr_id_commit[1].rs1 ;
  wire [5:0] \commit_instr_id_commit[1].rs1_t0 ;
  wire [5:0] \commit_instr_id_commit[1].rs1_t1 ;
  wire [5:0] \commit_instr_id_commit[1].rs2 ;
  wire [5:0] \commit_instr_id_commit[1].rs2_t0 ;
  wire [5:0] \commit_instr_id_commit[1].rs2_t1 ;
  wire [1:0] \commit_instr_id_commit[1].trans_id ;
  wire [1:0] \commit_instr_id_commit[1].trans_id_t0 ;
  wire [1:0] \commit_instr_id_commit[1].trans_id_t1 ;
  wire \commit_instr_id_commit[1].use_imm ;
  wire \commit_instr_id_commit[1].use_imm_t0 ;
  wire \commit_instr_id_commit[1].use_imm_t1 ;
  wire \commit_instr_id_commit[1].use_pc ;
  wire \commit_instr_id_commit[1].use_pc_t0 ;
  wire \commit_instr_id_commit[1].use_pc_t1 ;
  wire \commit_instr_id_commit[1].use_zimm ;
  wire \commit_instr_id_commit[1].use_zimm_t0 ;
  wire \commit_instr_id_commit[1].use_zimm_t1 ;
  wire \commit_instr_id_commit[1].valid ;
  wire \commit_instr_id_commit[1].valid_t0 ;
  wire \commit_instr_id_commit[1].valid_t1 ;
  wire [11:0] csr_addr_ex_csr;
  wire [11:0] csr_addr_ex_csr_t0;
  wire [11:0] csr_addr_ex_csr_t1;
  wire csr_commit_commit_ex;
  wire csr_commit_commit_ex_t0;
  wire csr_commit_commit_ex_t1;
  wire [63:0] \csr_exception_csr_commit.cause ;
  wire [63:0] \csr_exception_csr_commit.cause_t0 ;
  wire [63:0] \csr_exception_csr_commit.cause_t1 ;
  wire [63:0] \csr_exception_csr_commit.tval ;
  wire [63:0] \csr_exception_csr_commit.tval_t0 ;
  wire [63:0] \csr_exception_csr_commit.tval_t1 ;
  wire \csr_exception_csr_commit.valid ;
  wire \csr_exception_csr_commit.valid_t0 ;
  wire \csr_exception_csr_commit.valid_t1 ;
  wire [6:0] csr_op_commit_csr;
  wire [6:0] csr_op_commit_csr_t0;
  wire [6:0] csr_op_commit_csr_t1;
  wire [63:0] csr_rdata_csr_commit;
  wire [63:0] csr_rdata_csr_commit_t0;
  wire [63:0] csr_rdata_csr_commit_t1;
  wire csr_valid_id_ex;
  wire csr_valid_id_ex_t0;
  wire csr_valid_id_ex_t1;
  wire [63:0] csr_wdata_commit_csr;
  wire [63:0] csr_wdata_commit_csr_t0;
  wire [63:0] csr_wdata_commit_csr_t1;
  wire csr_write_fflags_commit_cs;
  wire csr_write_fflags_commit_cs_t0;
  wire csr_write_fflags_commit_cs_t1;
  wire dcache_en_csr_nbdcache;
  wire dcache_en_csr_nbdcache_t0;
  wire dcache_en_csr_nbdcache_t1;
  wire dcache_flush_ack_cache_ctrl;
  wire dcache_flush_ack_cache_ctrl_t0;
  wire dcache_flush_ack_cache_ctrl_t1;
  wire dcache_flush_ctrl_cache;
  wire dcache_flush_ctrl_cache_t0;
  wire dcache_flush_ctrl_cache_t1;
  wire debug_mode;
  wire debug_mode_t0;
  wire debug_mode_t1;
  wire debug_req_i;
  wire debug_req_i_t0;
  wire debug_req_i_t1;
  wire dirty_fp_state;
  wire dirty_fp_state_t0;
  wire dirty_fp_state_t1;
  wire en_ld_st_translation_csr_ex;
  wire en_ld_st_translation_csr_ex_t0;
  wire en_ld_st_translation_csr_ex_t1;
  wire enable_translation_csr_ex;
  wire enable_translation_csr_ex_t0;
  wire enable_translation_csr_ex_t1;
  wire [63:0] epc_commit_pcgen;
  wire [63:0] epc_commit_pcgen_t0;
  wire [63:0] epc_commit_pcgen_t1;
  wire eret;
  wire eret_t0;
  wire eret_t1;
  wire [63:0] \ex_commit.cause ;
  wire [63:0] \ex_commit.cause_t0 ;
  wire [63:0] \ex_commit.cause_t1 ;
  wire [63:0] \ex_commit.tval ;
  wire [63:0] \ex_commit.tval_t0 ;
  wire [63:0] \ex_commit.tval_t1 ;
  wire \ex_commit.valid ;
  wire \ex_commit.valid_t0 ;
  wire \ex_commit.valid_t1 ;
  wire fence_commit_controller;
  wire fence_commit_controller_t0;
  wire fence_commit_controller_t1;
  wire fence_i_commit_controller;
  wire fence_i_commit_controller_t0;
  wire fence_i_commit_controller_t1;
  wire [63:0] \fetch_entry_if_id.address ;
  wire [63:0] \fetch_entry_if_id.address_t0 ;
  wire [63:0] \fetch_entry_if_id.address_t1 ;
  wire [2:0] \fetch_entry_if_id.branch_predict.cf ;
  wire [2:0] \fetch_entry_if_id.branch_predict.cf_t0 ;
  wire [2:0] \fetch_entry_if_id.branch_predict.cf_t1 ;
  wire [63:0] \fetch_entry_if_id.branch_predict.predict_address ;
  wire [63:0] \fetch_entry_if_id.branch_predict.predict_address_t0 ;
  wire [63:0] \fetch_entry_if_id.branch_predict.predict_address_t1 ;
  wire [63:0] \fetch_entry_if_id.ex.cause ;
  wire [63:0] \fetch_entry_if_id.ex.cause_t0 ;
  wire [63:0] \fetch_entry_if_id.ex.cause_t1 ;
  wire [63:0] \fetch_entry_if_id.ex.tval ;
  wire [63:0] \fetch_entry_if_id.ex.tval_t0 ;
  wire [63:0] \fetch_entry_if_id.ex.tval_t1 ;
  wire \fetch_entry_if_id.ex.valid ;
  wire \fetch_entry_if_id.ex.valid_t0 ;
  wire \fetch_entry_if_id.ex.valid_t1 ;
  wire [31:0] \fetch_entry_if_id.instruction ;
  wire [31:0] \fetch_entry_if_id.instruction_t0 ;
  wire [31:0] \fetch_entry_if_id.instruction_t1 ;
  wire fetch_ready_id_if;
  wire fetch_ready_id_if_t0;
  wire fetch_ready_id_if_t1;
  wire fetch_valid_if_id;
  wire fetch_valid_if_id_t0;
  wire fetch_valid_if_id_t1;
  wire [4:0] fflags_csr_commit;
  wire [4:0] fflags_csr_commit_t0;
  wire [4:0] fflags_csr_commit_t1;
  wire [63:0] \flu_exception_ex_id.cause ;
  wire [63:0] \flu_exception_ex_id.cause_t0 ;
  wire [63:0] \flu_exception_ex_id.cause_t1 ;
  wire [63:0] \flu_exception_ex_id.tval ;
  wire [63:0] \flu_exception_ex_id.tval_t0 ;
  wire [63:0] \flu_exception_ex_id.tval_t1 ;
  wire \flu_exception_ex_id.valid ;
  wire \flu_exception_ex_id.valid_t0 ;
  wire \flu_exception_ex_id.valid_t1 ;
  wire flu_ready_ex_id;
  wire flu_ready_ex_id_t0;
  wire flu_ready_ex_id_t1;
  wire [63:0] flu_result_ex_id;
  wire [63:0] flu_result_ex_id_t0;
  wire [63:0] flu_result_ex_id_t1;
  wire [1:0] flu_trans_id_ex_id;
  wire [1:0] flu_trans_id_ex_id_t0;
  wire [1:0] flu_trans_id_ex_id_t1;
  wire flu_valid_ex_id;
  wire flu_valid_ex_id_t0;
  wire flu_valid_ex_id_t1;
  wire flush_commit;
  wire flush_commit_t0;
  wire flush_commit_t1;
  wire flush_csr_ctrl;
  wire flush_csr_ctrl_t0;
  wire flush_csr_ctrl_t1;
  wire flush_ctrl_bp;
  wire flush_ctrl_bp_t0;
  wire flush_ctrl_bp_t1;
  wire flush_ctrl_ex;
  wire flush_ctrl_ex_t0;
  wire flush_ctrl_ex_t1;
  wire flush_ctrl_id;
  wire flush_ctrl_id_t0;
  wire flush_ctrl_id_t1;
  wire flush_ctrl_if;
  wire flush_ctrl_if_t0;
  wire flush_ctrl_if_t1;
  wire flush_tlb_ctrl_ex;
  wire flush_tlb_ctrl_ex_t0;
  wire flush_tlb_ctrl_ex_t1;
  wire flush_unissued_instr_ctrl_id;
  wire flush_unissued_instr_ctrl_id_t0;
  wire flush_unissued_instr_ctrl_id_t1;
  wire [6:0] fprec_csr_ex;
  wire [6:0] fprec_csr_ex_t0;
  wire [6:0] fprec_csr_ex_t1;
  wire [63:0] \fpu_exception_ex_id.cause ;
  wire [63:0] \fpu_exception_ex_id.cause_t0 ;
  wire [63:0] \fpu_exception_ex_id.cause_t1 ;
  wire [63:0] \fpu_exception_ex_id.tval ;
  wire [63:0] \fpu_exception_ex_id.tval_t0 ;
  wire [63:0] \fpu_exception_ex_id.tval_t1 ;
  wire \fpu_exception_ex_id.valid ;
  wire \fpu_exception_ex_id.valid_t0 ;
  wire \fpu_exception_ex_id.valid_t1 ;
  wire [1:0] fpu_fmt_id_ex;
  wire [1:0] fpu_fmt_id_ex_t0;
  wire [1:0] fpu_fmt_id_ex_t1;
  wire fpu_ready_ex_id;
  wire fpu_ready_ex_id_t0;
  wire fpu_ready_ex_id_t1;
  wire [63:0] fpu_result_ex_id;
  wire [63:0] fpu_result_ex_id_t0;
  wire [63:0] fpu_result_ex_id_t1;
  wire [2:0] fpu_rm_id_ex;
  wire [2:0] fpu_rm_id_ex_t0;
  wire [2:0] fpu_rm_id_ex_t1;
  wire [1:0] fpu_trans_id_ex_id;
  wire [1:0] fpu_trans_id_ex_id_t0;
  wire [1:0] fpu_trans_id_ex_id_t1;
  wire fpu_valid_ex_id;
  wire fpu_valid_ex_id_t0;
  wire fpu_valid_ex_id_t1;
  wire fpu_valid_id_ex;
  wire fpu_valid_id_ex_t0;
  wire fpu_valid_id_ex_t1;
  wire [2:0] frm_csr_id_issue_ex;
  wire [2:0] frm_csr_id_issue_ex_t0;
  wire [2:0] frm_csr_id_issue_ex_t1;
  wire [1:0] fs;
  wire [1:0] fs_t0;
  wire [1:0] fs_t1;
  wire [3:0] \fu_data_id_ex.fu ;
  wire [3:0] \fu_data_id_ex.fu_t0 ;
  wire [3:0] \fu_data_id_ex.fu_t1 ;
  wire [63:0] \fu_data_id_ex.imm ;
  wire [63:0] \fu_data_id_ex.imm_t0 ;
  wire [63:0] \fu_data_id_ex.imm_t1 ;
  wire [63:0] \fu_data_id_ex.operand_a ;
  wire [63:0] \fu_data_id_ex.operand_a_t0 ;
  wire [63:0] \fu_data_id_ex.operand_a_t1 ;
  wire [63:0] \fu_data_id_ex.operand_b ;
  wire [63:0] \fu_data_id_ex.operand_b_t0 ;
  wire [63:0] \fu_data_id_ex.operand_b_t1 ;
  wire [6:0] \fu_data_id_ex.operator ;
  wire [6:0] \fu_data_id_ex.operator_t0 ;
  wire [6:0] \fu_data_id_ex.operator_t1 ;
  wire [1:0] \fu_data_id_ex.trans_id ;
  wire [1:0] \fu_data_id_ex.trans_id_t0 ;
  wire [1:0] \fu_data_id_ex.trans_id_t1 ;
  wire halt_csr_ctrl;
  wire halt_csr_ctrl_t0;
  wire halt_csr_ctrl_t1;
  wire halt_ctrl;
  wire halt_ctrl_t0;
  wire halt_ctrl_t1;
  wire [63:0] hart_id_i;
  wire [63:0] hart_id_i_t0;
  wire [63:0] hart_id_i_t1;
  wire icache_en_csr;
  wire icache_en_csr_t0;
  wire icache_en_csr_t1;
  wire icache_flush_ctrl_cache;
  wire icache_flush_ctrl_cache_t0;
  wire icache_flush_ctrl_cache_t1;
  wire ipi_i;
  wire ipi_i_t0;
  wire ipi_i_t1;
  wire \irq_ctrl_csr_id.global_enable ;
  wire \irq_ctrl_csr_id.global_enable_t0 ;
  wire \irq_ctrl_csr_id.global_enable_t1 ;
  wire [63:0] \irq_ctrl_csr_id.mideleg ;
  wire [63:0] \irq_ctrl_csr_id.mideleg_t0 ;
  wire [63:0] \irq_ctrl_csr_id.mideleg_t1 ;
  wire [63:0] \irq_ctrl_csr_id.mie ;
  wire [63:0] \irq_ctrl_csr_id.mie_t0 ;
  wire [63:0] \irq_ctrl_csr_id.mie_t1 ;
  wire [63:0] \irq_ctrl_csr_id.mip ;
  wire [63:0] \irq_ctrl_csr_id.mip_t0 ;
  wire [63:0] \irq_ctrl_csr_id.mip_t1 ;
  wire \irq_ctrl_csr_id.sie ;
  wire \irq_ctrl_csr_id.sie_t0 ;
  wire \irq_ctrl_csr_id.sie_t1 ;
  wire [1:0] irq_i;
  wire [1:0] irq_i_t0;
  wire [1:0] irq_i_t1;
  wire is_compressed_instr_id_ex;
  wire is_compressed_instr_id_ex_t0;
  wire is_compressed_instr_id_ex_t1;
  wire is_ctrl_fow_id_issue;
  wire is_ctrl_fow_id_issue_t0;
  wire is_ctrl_fow_id_issue_t1;
  wire [2:0] \issue_entry_id_issue.bp.cf ;
  wire [2:0] \issue_entry_id_issue.bp.cf_t0 ;
  wire [2:0] \issue_entry_id_issue.bp.cf_t1 ;
  wire [63:0] \issue_entry_id_issue.bp.predict_address ;
  wire [63:0] \issue_entry_id_issue.bp.predict_address_t0 ;
  wire [63:0] \issue_entry_id_issue.bp.predict_address_t1 ;
  wire [63:0] \issue_entry_id_issue.ex.cause ;
  wire [63:0] \issue_entry_id_issue.ex.cause_t0 ;
  wire [63:0] \issue_entry_id_issue.ex.cause_t1 ;
  wire [63:0] \issue_entry_id_issue.ex.tval ;
  wire [63:0] \issue_entry_id_issue.ex.tval_t0 ;
  wire [63:0] \issue_entry_id_issue.ex.tval_t1 ;
  wire \issue_entry_id_issue.ex.valid ;
  wire \issue_entry_id_issue.ex.valid_t0 ;
  wire \issue_entry_id_issue.ex.valid_t1 ;
  wire [3:0] \issue_entry_id_issue.fu ;
  wire [3:0] \issue_entry_id_issue.fu_t0 ;
  wire [3:0] \issue_entry_id_issue.fu_t1 ;
  wire \issue_entry_id_issue.is_compressed ;
  wire \issue_entry_id_issue.is_compressed_t0 ;
  wire \issue_entry_id_issue.is_compressed_t1 ;
  wire [6:0] \issue_entry_id_issue.op ;
  wire [6:0] \issue_entry_id_issue.op_t0 ;
  wire [6:0] \issue_entry_id_issue.op_t1 ;
  wire [63:0] \issue_entry_id_issue.pc ;
  wire [63:0] \issue_entry_id_issue.pc_t0 ;
  wire [63:0] \issue_entry_id_issue.pc_t1 ;
  wire [5:0] \issue_entry_id_issue.rd ;
  wire [5:0] \issue_entry_id_issue.rd_t0 ;
  wire [5:0] \issue_entry_id_issue.rd_t1 ;
  wire [63:0] \issue_entry_id_issue.result ;
  wire [63:0] \issue_entry_id_issue.result_t0 ;
  wire [63:0] \issue_entry_id_issue.result_t1 ;
  wire [5:0] \issue_entry_id_issue.rs1 ;
  wire [5:0] \issue_entry_id_issue.rs1_t0 ;
  wire [5:0] \issue_entry_id_issue.rs1_t1 ;
  wire [5:0] \issue_entry_id_issue.rs2 ;
  wire [5:0] \issue_entry_id_issue.rs2_t0 ;
  wire [5:0] \issue_entry_id_issue.rs2_t1 ;
  wire [1:0] \issue_entry_id_issue.trans_id ;
  wire [1:0] \issue_entry_id_issue.trans_id_t0 ;
  wire [1:0] \issue_entry_id_issue.trans_id_t1 ;
  wire \issue_entry_id_issue.use_imm ;
  wire \issue_entry_id_issue.use_imm_t0 ;
  wire \issue_entry_id_issue.use_imm_t1 ;
  wire \issue_entry_id_issue.use_pc ;
  wire \issue_entry_id_issue.use_pc_t0 ;
  wire \issue_entry_id_issue.use_pc_t1 ;
  wire \issue_entry_id_issue.use_zimm ;
  wire \issue_entry_id_issue.use_zimm_t0 ;
  wire \issue_entry_id_issue.use_zimm_t1 ;
  wire \issue_entry_id_issue.valid ;
  wire \issue_entry_id_issue.valid_t0 ;
  wire \issue_entry_id_issue.valid_t1 ;
  wire issue_entry_valid_id_issue;
  wire issue_entry_valid_id_issue_t0;
  wire issue_entry_valid_id_issue_t1;
  wire issue_instr_issue_id;
  wire issue_instr_issue_id_t0;
  wire issue_instr_issue_id_t1;
  wire [1:0] ld_st_priv_lvl_csr_ex;
  wire [1:0] ld_st_priv_lvl_csr_ex_t0;
  wire [1:0] ld_st_priv_lvl_csr_ex_t1;
  wire [63:0] \load_exception_ex_id.cause ;
  wire [63:0] \load_exception_ex_id.cause_t0 ;
  wire [63:0] \load_exception_ex_id.cause_t1 ;
  wire [63:0] \load_exception_ex_id.tval ;
  wire [63:0] \load_exception_ex_id.tval_t0 ;
  wire [63:0] \load_exception_ex_id.tval_t1 ;
  wire \load_exception_ex_id.valid ;
  wire \load_exception_ex_id.valid_t0 ;
  wire \load_exception_ex_id.valid_t1 ;
  wire [63:0] load_result_ex_id;
  wire [63:0] load_result_ex_id_t0;
  wire [63:0] load_result_ex_id_t1;
  wire [1:0] load_trans_id_ex_id;
  wire [1:0] load_trans_id_ex_id_t0;
  wire [1:0] load_trans_id_ex_id_t1;
  wire load_valid_ex_id;
  wire load_valid_ex_id_t0;
  wire load_valid_ex_id_t1;
  wire lsu_commit_commit_ex;
  wire lsu_commit_commit_ex_t0;
  wire lsu_commit_commit_ex_t1;
  wire lsu_commit_ready_ex_commit;
  wire lsu_commit_ready_ex_commit_t0;
  wire lsu_commit_ready_ex_commit_t1;
  wire [1:0] lsu_commit_trans_id;
  wire [1:0] lsu_commit_trans_id_t0;
  wire [1:0] lsu_commit_trans_id_t1;
  wire lsu_ready_ex_id;
  wire lsu_ready_ex_id_t0;
  wire lsu_ready_ex_id_t1;
  wire lsu_valid_id_ex;
  wire lsu_valid_id_ex_t0;
  wire lsu_valid_id_ex_t1;
  wire mult_valid_id_ex;
  wire mult_valid_id_ex_t0;
  wire mult_valid_id_ex_t1;
  wire mxr_csr_ex;
  wire mxr_csr_ex_t0;
  wire mxr_csr_ex_t1;
  wire no_st_pending_commit;
  wire no_st_pending_commit_t0;
  wire no_st_pending_commit_t1;
  wire no_st_pending_ex;
  wire no_st_pending_ex_t0;
  wire no_st_pending_ex_t1;
  wire [63:0] pc_commit;
  wire [63:0] pc_commit_t0;
  wire [63:0] pc_commit_t1;
  wire [63:0] pc_id_ex;
  wire [63:0] pc_id_ex_t0;
  wire [63:0] pc_id_ex_t1;
  wire [1:0] priv_lvl;
  wire [1:0] priv_lvl_t0;
  wire [1:0] priv_lvl_t1;
  wire [31:0] read_instr;
  wire resolve_branch_ex_id;
  wire resolve_branch_ex_id_t0;
  wire resolve_branch_ex_id_t1;
  wire [2:0] \resolved_branch.cf_type ;
  wire [2:0] \resolved_branch.cf_type_t0 ;
  wire [2:0] \resolved_branch.cf_type_t1 ;
  wire \resolved_branch.is_mispredict ;
  wire \resolved_branch.is_mispredict_t0 ;
  wire \resolved_branch.is_mispredict_t1 ;
  wire \resolved_branch.is_taken ;
  wire \resolved_branch.is_taken_t0 ;
  wire \resolved_branch.is_taken_t1 ;
  wire [63:0] \resolved_branch.pc ;
  wire [63:0] \resolved_branch.pc_t0 ;
  wire [63:0] \resolved_branch.pc_t1 ;
  wire [63:0] \resolved_branch.target_address ;
  wire [63:0] \resolved_branch.target_address_t0 ;
  wire [63:0] \resolved_branch.target_address_t1 ;
  wire \resolved_branch.valid ;
  wire \resolved_branch.valid_t0 ;
  wire \resolved_branch.valid_t1 ;
  wire [63:0] rs1_forwarding_id_ex;
  wire [63:0] rs1_forwarding_id_ex_t0;
  wire [63:0] rs1_forwarding_id_ex_t1;
  wire [63:0] rs2_forwarding_id_ex;
  wire [63:0] rs2_forwarding_id_ex_t0;
  wire [63:0] rs2_forwarding_id_ex_t1;
  wire [43:0] satp_ppn_csr_ex;
  wire [43:0] satp_ppn_csr_ex_t0;
  wire [43:0] satp_ppn_csr_ex_t1;
  wire sb_full;
  wire sb_full_t0;
  wire sb_full_t1;
  wire set_debug_pc;
  wire set_debug_pc_t0;
  wire set_debug_pc_t1;
  wire set_pc_ctrl_pcgen;
  wire set_pc_ctrl_pcgen_t0;
  wire set_pc_ctrl_pcgen_t1;
  wire sfence_vma_commit_controller;
  wire sfence_vma_commit_controller_t0;
  wire sfence_vma_commit_controller_t1;
  wire single_step_csr_commit;
  wire single_step_csr_commit_t0;
  wire single_step_csr_commit_t1;
  wire [63:0] \store_exception_ex_id.cause ;
  wire [63:0] \store_exception_ex_id.cause_t0 ;
  wire [63:0] \store_exception_ex_id.cause_t1 ;
  wire [63:0] \store_exception_ex_id.tval ;
  wire [63:0] \store_exception_ex_id.tval_t0 ;
  wire [63:0] \store_exception_ex_id.tval_t1 ;
  wire \store_exception_ex_id.valid ;
  wire \store_exception_ex_id.valid_t0 ;
  wire \store_exception_ex_id.valid_t1 ;
  wire [63:0] store_result_ex_id;
  wire [63:0] store_result_ex_id_t0;
  wire [63:0] store_result_ex_id_t1;
  wire [1:0] store_trans_id_ex_id;
  wire [1:0] store_trans_id_ex_id_t0;
  wire [1:0] store_trans_id_ex_id_t1;
  wire store_valid_ex_id;
  wire store_valid_ex_id_t0;
  wire store_valid_ex_id_t1;
  wire sum_csr_ex;
  wire sum_csr_ex_t0;
  wire sum_csr_ex_t1;
  wire time_irq_i;
  wire time_irq_i_t0;
  wire time_irq_i_t1;
  wire [31:0] \tmp_icache_dreq_cache_if.data ;
  wire [31:0] \tmp_icache_dreq_cache_if.data_t0 ;
  wire [31:0] \tmp_icache_dreq_cache_if.data_t1 ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.cause ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.cause_t0 ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.cause_t1 ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.tval ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.tval_t0 ;
  wire [63:0] \tmp_icache_dreq_cache_if.ex.tval_t1 ;
  wire \tmp_icache_dreq_cache_if.ex.valid ;
  wire \tmp_icache_dreq_cache_if.ex.valid_t0 ;
  wire \tmp_icache_dreq_cache_if.ex.valid_t1 ;
  wire \tmp_icache_dreq_cache_if.ready ;
  wire \tmp_icache_dreq_cache_if.ready_t0 ;
  wire \tmp_icache_dreq_cache_if.ready_t1 ;
  wire [63:0] \tmp_icache_dreq_cache_if.vaddr ;
  wire [63:0] \tmp_icache_dreq_cache_if.vaddr_t0 ;
  wire [63:0] \tmp_icache_dreq_cache_if.vaddr_t1 ;
  wire \tmp_icache_dreq_cache_if.valid ;
  wire \tmp_icache_dreq_cache_if.valid_t0 ;
  wire \tmp_icache_dreq_cache_if.valid_t1 ;
  wire \tmp_icache_dreq_if_cache.kill_s1 ;
  wire \tmp_icache_dreq_if_cache.kill_s1_t0 ;
  wire \tmp_icache_dreq_if_cache.kill_s1_t1 ;
  wire \tmp_icache_dreq_if_cache.kill_s2 ;
  wire \tmp_icache_dreq_if_cache.kill_s2_t0 ;
  wire \tmp_icache_dreq_if_cache.kill_s2_t1 ;
  wire \tmp_icache_dreq_if_cache.req ;
  wire \tmp_icache_dreq_if_cache.req_t0 ;
  wire \tmp_icache_dreq_if_cache.req_t1 ;
  wire \tmp_icache_dreq_if_cache.spec ;
  wire \tmp_icache_dreq_if_cache.spec_t0 ;
  wire \tmp_icache_dreq_if_cache.spec_t1 ;
  wire [63:0] \tmp_icache_dreq_if_cache.vaddr ;
  wire [63:0] \tmp_icache_dreq_if_cache.vaddr_t0 ;
  wire [63:0] \tmp_icache_dreq_if_cache.vaddr_t1 ;
  wire [63:0] trap_vector_base_commit_pcgen;
  wire [63:0] trap_vector_base_commit_pcgen_t0;
  wire [63:0] trap_vector_base_commit_pcgen_t1;
  wire tsr_csr_id;
  wire tsr_csr_id_t0;
  wire tsr_csr_id_t1;
  wire tvm_csr_id;
  wire tvm_csr_id_t0;
  wire tvm_csr_id_t1;
  wire tw_csr_id;
  wire tw_csr_id_t0;
  wire tw_csr_id_t1;
  wire [4:0] \waddr_commit_id[0] ;
  wire [4:0] \waddr_commit_id[0]_t0 ;
  wire [4:0] \waddr_commit_id[0]_t1 ;
  wire [4:0] \waddr_commit_id[1] ;
  wire [4:0] \waddr_commit_id[1]_t0 ;
  wire [4:0] \waddr_commit_id[1]_t1 ;
  wire [63:0] \wdata_commit_id[0] ;
  wire [63:0] \wdata_commit_id[0]_t0 ;
  wire [63:0] \wdata_commit_id[0]_t1 ;
  wire [63:0] \wdata_commit_id[1] ;
  wire [63:0] \wdata_commit_id[1]_t0 ;
  wire [63:0] \wdata_commit_id[1]_t1 ;
  wire [1:0] we_fpr_commit_id;
  wire [1:0] we_fpr_commit_id_t0;
  wire [1:0] we_fpr_commit_id_t1;
  wire [1:0] we_gpr_commit_id;
  wire [1:0] we_gpr_commit_id_t0;
  wire [1:0] we_gpr_commit_id_t1;
  reg [4:0] prev_req [0:0];
  reg [255:0] prev_vaddr [0:0];
  assign dcache_flush_ack_cache_ctrl = 1'h1; // _BUF_, assign Y = A
  assign no_st_pending_commit = no_st_pending_ex; // _BUF_, assign Y = A
  assign debug_req_i = 1'h0; // _BUF_, assign Y = A
  assign time_irq_i = 1'h0; // _BUF_, assign Y = A
  assign ipi_i = 1'h0; // _BUF_, assign Y = A
  \commit_stage(NR_COMMIT_PORTS=32'b010)  commit_stage_i (
    .\amo_resp_i.ack (\amo_resp.ack ),
    .\amo_resp_i.ack_t0 (\amo_resp.ack_t0 ),
    .\amo_resp_i.ack_t1 (\amo_resp.ack_t1 ),
    .\amo_resp_i.result (\amo_resp.result ),
    .\amo_resp_i.result_t0 (\amo_resp.result_t0 ),
    .\amo_resp_i.result_t1 (\amo_resp.result_t1 ),
    .amo_valid_commit_o(amo_valid_commit),
    .amo_valid_commit_o_t0(amo_valid_commit_t0),
    .amo_valid_commit_o_t1(amo_valid_commit_t1),
    .clk_i(clk_i),
    .commit_ack_o(commit_ack),
    .commit_ack_o_t0(commit_ack_t0),
    .commit_ack_o_t1(commit_ack_t1),
    .commit_csr_o(csr_commit_commit_ex),
    .commit_csr_o_t0(csr_commit_commit_ex_t0),
    .commit_csr_o_t1(csr_commit_commit_ex_t1),
    .\commit_instr_i[0].bp.cf (\commit_instr_id_commit[0].bp.cf ),
    .\commit_instr_i[0].bp.cf_t0 (\commit_instr_id_commit[0].bp.cf_t0 ),
    .\commit_instr_i[0].bp.cf_t1 (\commit_instr_id_commit[0].bp.cf_t1 ),
    .\commit_instr_i[0].bp.predict_address (\commit_instr_id_commit[0].bp.predict_address ),
    .\commit_instr_i[0].bp.predict_address_t0 (\commit_instr_id_commit[0].bp.predict_address_t0 ),
    .\commit_instr_i[0].bp.predict_address_t1 (\commit_instr_id_commit[0].bp.predict_address_t1 ),
    .\commit_instr_i[0].ex.cause (\commit_instr_id_commit[0].ex.cause ),
    .\commit_instr_i[0].ex.cause_t0 (\commit_instr_id_commit[0].ex.cause_t0 ),
    .\commit_instr_i[0].ex.cause_t1 (\commit_instr_id_commit[0].ex.cause_t1 ),
    .\commit_instr_i[0].ex.tval (\commit_instr_id_commit[0].ex.tval ),
    .\commit_instr_i[0].ex.tval_t0 (\commit_instr_id_commit[0].ex.tval_t0 ),
    .\commit_instr_i[0].ex.tval_t1 (\commit_instr_id_commit[0].ex.tval_t1 ),
    .\commit_instr_i[0].ex.valid (\commit_instr_id_commit[0].ex.valid ),
    .\commit_instr_i[0].ex.valid_t0 (\commit_instr_id_commit[0].ex.valid_t0 ),
    .\commit_instr_i[0].ex.valid_t1 (\commit_instr_id_commit[0].ex.valid_t1 ),
    .\commit_instr_i[0].fu (\commit_instr_id_commit[0].fu ),
    .\commit_instr_i[0].fu_t0 (\commit_instr_id_commit[0].fu_t0 ),
    .\commit_instr_i[0].fu_t1 (\commit_instr_id_commit[0].fu_t1 ),
    .\commit_instr_i[0].is_compressed (\commit_instr_id_commit[0].is_compressed ),
    .\commit_instr_i[0].is_compressed_t0 (\commit_instr_id_commit[0].is_compressed_t0 ),
    .\commit_instr_i[0].is_compressed_t1 (\commit_instr_id_commit[0].is_compressed_t1 ),
    .\commit_instr_i[0].op (\commit_instr_id_commit[0].op ),
    .\commit_instr_i[0].op_t0 (\commit_instr_id_commit[0].op_t0 ),
    .\commit_instr_i[0].op_t1 (\commit_instr_id_commit[0].op_t1 ),
    .\commit_instr_i[0].pc (\commit_instr_id_commit[0].pc ),
    .\commit_instr_i[0].pc_t0 (\commit_instr_id_commit[0].pc_t0 ),
    .\commit_instr_i[0].pc_t1 (\commit_instr_id_commit[0].pc_t1 ),
    .\commit_instr_i[0].rd (\commit_instr_id_commit[0].rd ),
    .\commit_instr_i[0].rd_t0 (\commit_instr_id_commit[0].rd_t0 ),
    .\commit_instr_i[0].rd_t1 (\commit_instr_id_commit[0].rd_t1 ),
    .\commit_instr_i[0].result (\commit_instr_id_commit[0].result ),
    .\commit_instr_i[0].result_t0 (\commit_instr_id_commit[0].result_t0 ),
    .\commit_instr_i[0].result_t1 (\commit_instr_id_commit[0].result_t1 ),
    .\commit_instr_i[0].rs1 (\commit_instr_id_commit[0].rs1 ),
    .\commit_instr_i[0].rs1_t0 (\commit_instr_id_commit[0].rs1_t0 ),
    .\commit_instr_i[0].rs1_t1 (\commit_instr_id_commit[0].rs1_t1 ),
    .\commit_instr_i[0].rs2 (\commit_instr_id_commit[0].rs2 ),
    .\commit_instr_i[0].rs2_t0 (\commit_instr_id_commit[0].rs2_t0 ),
    .\commit_instr_i[0].rs2_t1 (\commit_instr_id_commit[0].rs2_t1 ),
    .\commit_instr_i[0].trans_id (\commit_instr_id_commit[0].trans_id ),
    .\commit_instr_i[0].trans_id_t0 (\commit_instr_id_commit[0].trans_id_t0 ),
    .\commit_instr_i[0].trans_id_t1 (\commit_instr_id_commit[0].trans_id_t1 ),
    .\commit_instr_i[0].use_imm (\commit_instr_id_commit[0].use_imm ),
    .\commit_instr_i[0].use_imm_t0 (\commit_instr_id_commit[0].use_imm_t0 ),
    .\commit_instr_i[0].use_imm_t1 (\commit_instr_id_commit[0].use_imm_t1 ),
    .\commit_instr_i[0].use_pc (\commit_instr_id_commit[0].use_pc ),
    .\commit_instr_i[0].use_pc_t0 (\commit_instr_id_commit[0].use_pc_t0 ),
    .\commit_instr_i[0].use_pc_t1 (\commit_instr_id_commit[0].use_pc_t1 ),
    .\commit_instr_i[0].use_zimm (\commit_instr_id_commit[0].use_zimm ),
    .\commit_instr_i[0].use_zimm_t0 (\commit_instr_id_commit[0].use_zimm_t0 ),
    .\commit_instr_i[0].use_zimm_t1 (\commit_instr_id_commit[0].use_zimm_t1 ),
    .\commit_instr_i[0].valid (\commit_instr_id_commit[0].valid ),
    .\commit_instr_i[0].valid_t0 (\commit_instr_id_commit[0].valid_t0 ),
    .\commit_instr_i[0].valid_t1 (\commit_instr_id_commit[0].valid_t1 ),
    .\commit_instr_i[1].bp.cf (\commit_instr_id_commit[1].bp.cf ),
    .\commit_instr_i[1].bp.cf_t0 (\commit_instr_id_commit[1].bp.cf_t0 ),
    .\commit_instr_i[1].bp.cf_t1 (\commit_instr_id_commit[1].bp.cf_t1 ),
    .\commit_instr_i[1].bp.predict_address (\commit_instr_id_commit[1].bp.predict_address ),
    .\commit_instr_i[1].bp.predict_address_t0 (\commit_instr_id_commit[1].bp.predict_address_t0 ),
    .\commit_instr_i[1].bp.predict_address_t1 (\commit_instr_id_commit[1].bp.predict_address_t1 ),
    .\commit_instr_i[1].ex.cause (\commit_instr_id_commit[1].ex.cause ),
    .\commit_instr_i[1].ex.cause_t0 (\commit_instr_id_commit[1].ex.cause_t0 ),
    .\commit_instr_i[1].ex.cause_t1 (\commit_instr_id_commit[1].ex.cause_t1 ),
    .\commit_instr_i[1].ex.tval (\commit_instr_id_commit[1].ex.tval ),
    .\commit_instr_i[1].ex.tval_t0 (\commit_instr_id_commit[1].ex.tval_t0 ),
    .\commit_instr_i[1].ex.tval_t1 (\commit_instr_id_commit[1].ex.tval_t1 ),
    .\commit_instr_i[1].ex.valid (\commit_instr_id_commit[1].ex.valid ),
    .\commit_instr_i[1].ex.valid_t0 (\commit_instr_id_commit[1].ex.valid_t0 ),
    .\commit_instr_i[1].ex.valid_t1 (\commit_instr_id_commit[1].ex.valid_t1 ),
    .\commit_instr_i[1].fu (\commit_instr_id_commit[1].fu ),
    .\commit_instr_i[1].fu_t0 (\commit_instr_id_commit[1].fu_t0 ),
    .\commit_instr_i[1].fu_t1 (\commit_instr_id_commit[1].fu_t1 ),
    .\commit_instr_i[1].is_compressed (\commit_instr_id_commit[1].is_compressed ),
    .\commit_instr_i[1].is_compressed_t0 (\commit_instr_id_commit[1].is_compressed_t0 ),
    .\commit_instr_i[1].is_compressed_t1 (\commit_instr_id_commit[1].is_compressed_t1 ),
    .\commit_instr_i[1].op (\commit_instr_id_commit[1].op ),
    .\commit_instr_i[1].op_t0 (\commit_instr_id_commit[1].op_t0 ),
    .\commit_instr_i[1].op_t1 (\commit_instr_id_commit[1].op_t1 ),
    .\commit_instr_i[1].pc (\commit_instr_id_commit[1].pc ),
    .\commit_instr_i[1].pc_t0 (\commit_instr_id_commit[1].pc_t0 ),
    .\commit_instr_i[1].pc_t1 (\commit_instr_id_commit[1].pc_t1 ),
    .\commit_instr_i[1].rd (\commit_instr_id_commit[1].rd ),
    .\commit_instr_i[1].rd_t0 (\commit_instr_id_commit[1].rd_t0 ),
    .\commit_instr_i[1].rd_t1 (\commit_instr_id_commit[1].rd_t1 ),
    .\commit_instr_i[1].result (\commit_instr_id_commit[1].result ),
    .\commit_instr_i[1].result_t0 (\commit_instr_id_commit[1].result_t0 ),
    .\commit_instr_i[1].result_t1 (\commit_instr_id_commit[1].result_t1 ),
    .\commit_instr_i[1].rs1 (\commit_instr_id_commit[1].rs1 ),
    .\commit_instr_i[1].rs1_t0 (\commit_instr_id_commit[1].rs1_t0 ),
    .\commit_instr_i[1].rs1_t1 (\commit_instr_id_commit[1].rs1_t1 ),
    .\commit_instr_i[1].rs2 (\commit_instr_id_commit[1].rs2 ),
    .\commit_instr_i[1].rs2_t0 (\commit_instr_id_commit[1].rs2_t0 ),
    .\commit_instr_i[1].rs2_t1 (\commit_instr_id_commit[1].rs2_t1 ),
    .\commit_instr_i[1].trans_id (\commit_instr_id_commit[1].trans_id ),
    .\commit_instr_i[1].trans_id_t0 (\commit_instr_id_commit[1].trans_id_t0 ),
    .\commit_instr_i[1].trans_id_t1 (\commit_instr_id_commit[1].trans_id_t1 ),
    .\commit_instr_i[1].use_imm (\commit_instr_id_commit[1].use_imm ),
    .\commit_instr_i[1].use_imm_t0 (\commit_instr_id_commit[1].use_imm_t0 ),
    .\commit_instr_i[1].use_imm_t1 (\commit_instr_id_commit[1].use_imm_t1 ),
    .\commit_instr_i[1].use_pc (\commit_instr_id_commit[1].use_pc ),
    .\commit_instr_i[1].use_pc_t0 (\commit_instr_id_commit[1].use_pc_t0 ),
    .\commit_instr_i[1].use_pc_t1 (\commit_instr_id_commit[1].use_pc_t1 ),
    .\commit_instr_i[1].use_zimm (\commit_instr_id_commit[1].use_zimm ),
    .\commit_instr_i[1].use_zimm_t0 (\commit_instr_id_commit[1].use_zimm_t0 ),
    .\commit_instr_i[1].use_zimm_t1 (\commit_instr_id_commit[1].use_zimm_t1 ),
    .\commit_instr_i[1].valid (\commit_instr_id_commit[1].valid ),
    .\commit_instr_i[1].valid_t0 (\commit_instr_id_commit[1].valid_t0 ),
    .\commit_instr_i[1].valid_t1 (\commit_instr_id_commit[1].valid_t1 ),
    .commit_lsu_o(lsu_commit_commit_ex),
    .commit_lsu_o_t0(lsu_commit_commit_ex_t0),
    .commit_lsu_o_t1(lsu_commit_commit_ex_t1),
    .commit_lsu_ready_i(lsu_commit_ready_ex_commit),
    .commit_lsu_ready_i_t0(lsu_commit_ready_ex_commit_t0),
    .commit_lsu_ready_i_t1(lsu_commit_ready_ex_commit_t1),
    .commit_tran_id_o(lsu_commit_trans_id),
    .commit_tran_id_o_t0(lsu_commit_trans_id_t0),
    .commit_tran_id_o_t1(lsu_commit_trans_id_t1),
    .\csr_exception_i.cause (\csr_exception_csr_commit.cause ),
    .\csr_exception_i.cause_t0 (\csr_exception_csr_commit.cause_t0 ),
    .\csr_exception_i.cause_t1 (\csr_exception_csr_commit.cause_t1 ),
    .\csr_exception_i.tval (\csr_exception_csr_commit.tval ),
    .\csr_exception_i.tval_t0 (\csr_exception_csr_commit.tval_t0 ),
    .\csr_exception_i.tval_t1 (\csr_exception_csr_commit.tval_t1 ),
    .\csr_exception_i.valid (\csr_exception_csr_commit.valid ),
    .\csr_exception_i.valid_t0 (\csr_exception_csr_commit.valid_t0 ),
    .\csr_exception_i.valid_t1 (\csr_exception_csr_commit.valid_t1 ),
    .csr_op_o(csr_op_commit_csr),
    .csr_op_o_t0(csr_op_commit_csr_t0),
    .csr_op_o_t1(csr_op_commit_csr_t1),
    .csr_rdata_i(csr_rdata_csr_commit),
    .csr_rdata_i_t0(csr_rdata_csr_commit_t0),
    .csr_rdata_i_t1(csr_rdata_csr_commit_t1),
    .csr_wdata_o(csr_wdata_commit_csr),
    .csr_wdata_o_t0(csr_wdata_commit_csr_t0),
    .csr_wdata_o_t1(csr_wdata_commit_csr_t1),
    .csr_write_fflags_o(csr_write_fflags_commit_cs),
    .csr_write_fflags_o_t0(csr_write_fflags_commit_cs_t0),
    .csr_write_fflags_o_t1(csr_write_fflags_commit_cs_t1),
    .dirty_fp_state_o(dirty_fp_state),
    .dirty_fp_state_o_t0(dirty_fp_state_t0),
    .dirty_fp_state_o_t1(dirty_fp_state_t1),
    .\exception_o.cause (\ex_commit.cause ),
    .\exception_o.cause_t0 (\ex_commit.cause_t0 ),
    .\exception_o.cause_t1 (\ex_commit.cause_t1 ),
    .\exception_o.tval (\ex_commit.tval ),
    .\exception_o.tval_t0 (\ex_commit.tval_t0 ),
    .\exception_o.tval_t1 (\ex_commit.tval_t1 ),
    .\exception_o.valid (\ex_commit.valid ),
    .\exception_o.valid_t0 (\ex_commit.valid_t0 ),
    .\exception_o.valid_t1 (\ex_commit.valid_t1 ),
    .fence_i_o(fence_i_commit_controller),
    .fence_i_o_t0(fence_i_commit_controller_t0),
    .fence_i_o_t1(fence_i_commit_controller_t1),
    .fence_o(fence_commit_controller),
    .fence_o_t0(fence_commit_controller_t0),
    .fence_o_t1(fence_commit_controller_t1),
    .flush_commit_o(flush_commit),
    .flush_commit_o_t0(flush_commit_t0),
    .flush_commit_o_t1(flush_commit_t1),
    .flush_dcache_i(dcache_flush_ctrl_cache),
    .flush_dcache_i_t0(dcache_flush_ctrl_cache_t0),
    .flush_dcache_i_t1(dcache_flush_ctrl_cache_t1),
    .halt_i(halt_ctrl),
    .halt_i_t0(halt_ctrl_t0),
    .halt_i_t1(halt_ctrl_t1),
    .no_st_pending_i(no_st_pending_commit),
    .no_st_pending_i_t0(no_st_pending_commit_t0),
    .no_st_pending_i_t1(no_st_pending_commit_t1),
    .pc_o(pc_commit),
    .pc_o_t0(pc_commit_t0),
    .pc_o_t1(pc_commit_t1),
    .rst_ni(rst_ni),
    .sfence_vma_o(sfence_vma_commit_controller),
    .sfence_vma_o_t0(sfence_vma_commit_controller_t0),
    .sfence_vma_o_t1(sfence_vma_commit_controller_t1),
    .single_step_i(single_step_csr_commit),
    .single_step_i_t0(single_step_csr_commit_t0),
    .single_step_i_t1(single_step_csr_commit_t1),
    .\waddr_o[0] (\waddr_commit_id[0] ),
    .\waddr_o[0]_t0 (\waddr_commit_id[0]_t0 ),
    .\waddr_o[0]_t1 (\waddr_commit_id[0]_t1 ),
    .\waddr_o[1] (\waddr_commit_id[1] ),
    .\waddr_o[1]_t0 (\waddr_commit_id[1]_t0 ),
    .\waddr_o[1]_t1 (\waddr_commit_id[1]_t1 ),
    .\wdata_o[0] (\wdata_commit_id[0] ),
    .\wdata_o[0]_t0 (\wdata_commit_id[0]_t0 ),
    .\wdata_o[0]_t1 (\wdata_commit_id[0]_t1 ),
    .\wdata_o[1] (\wdata_commit_id[1] ),
    .\wdata_o[1]_t0 (\wdata_commit_id[1]_t0 ),
    .\wdata_o[1]_t1 (\wdata_commit_id[1]_t1 ),
    .we_fpr_o(we_fpr_commit_id),
    .we_fpr_o_t0(we_fpr_commit_id_t0),
    .we_fpr_o_t1(we_fpr_commit_id_t1),
    .we_gpr_o(we_gpr_commit_id),
    .we_gpr_o_t0(we_gpr_commit_id_t0),
    .we_gpr_o_t1(we_gpr_commit_id_t1)
  );
  controller controller_i (
    .clk_i(clk_i),
    .eret_i(eret),
    .eret_i_t0(eret_t0),
    .eret_i_t1(eret_t1),
    .ex_valid_i(\ex_commit.valid ),
    .ex_valid_i_t0(\ex_commit.valid_t0 ),
    .ex_valid_i_t1(\ex_commit.valid_t1 ),
    .fence_i(fence_commit_controller),
    .fence_i_i(fence_i_commit_controller),
    .fence_i_i_t0(fence_i_commit_controller_t0),
    .fence_i_i_t1(fence_i_commit_controller_t1),
    .fence_i_t0(fence_commit_controller_t0),
    .fence_i_t1(fence_commit_controller_t1),
    .flush_bp_o(flush_ctrl_bp),
    .flush_bp_o_t0(flush_ctrl_bp_t0),
    .flush_bp_o_t1(flush_ctrl_bp_t1),
    .flush_commit_i(flush_commit),
    .flush_commit_i_t0(flush_commit_t0),
    .flush_commit_i_t1(flush_commit_t1),
    .flush_csr_i(flush_csr_ctrl),
    .flush_csr_i_t0(flush_csr_ctrl_t0),
    .flush_csr_i_t1(flush_csr_ctrl_t1),
    .flush_dcache_ack_i(dcache_flush_ack_cache_ctrl),
    .flush_dcache_ack_i_t0(dcache_flush_ack_cache_ctrl_t0),
    .flush_dcache_ack_i_t1(dcache_flush_ack_cache_ctrl_t1),
    .flush_dcache_o(dcache_flush_ctrl_cache),
    .flush_dcache_o_t0(dcache_flush_ctrl_cache_t0),
    .flush_dcache_o_t1(dcache_flush_ctrl_cache_t1),
    .flush_ex_o(flush_ctrl_ex),
    .flush_ex_o_t0(flush_ctrl_ex_t0),
    .flush_ex_o_t1(flush_ctrl_ex_t1),
    .flush_icache_o(icache_flush_ctrl_cache),
    .flush_icache_o_t0(icache_flush_ctrl_cache_t0),
    .flush_icache_o_t1(icache_flush_ctrl_cache_t1),
    .flush_id_o(flush_ctrl_id),
    .flush_id_o_t0(flush_ctrl_id_t0),
    .flush_id_o_t1(flush_ctrl_id_t1),
    .flush_if_o(flush_ctrl_if),
    .flush_if_o_t0(flush_ctrl_if_t0),
    .flush_if_o_t1(flush_ctrl_if_t1),
    .flush_tlb_o(flush_tlb_ctrl_ex),
    .flush_tlb_o_t0(flush_tlb_ctrl_ex_t0),
    .flush_tlb_o_t1(flush_tlb_ctrl_ex_t1),
    .flush_unissued_instr_o(flush_unissued_instr_ctrl_id),
    .flush_unissued_instr_o_t0(flush_unissued_instr_ctrl_id_t0),
    .flush_unissued_instr_o_t1(flush_unissued_instr_ctrl_id_t1),
    .halt_csr_i(halt_csr_ctrl),
    .halt_csr_i_t0(halt_csr_ctrl_t0),
    .halt_csr_i_t1(halt_csr_ctrl_t1),
    .halt_o(halt_ctrl),
    .halt_o_t0(halt_ctrl_t0),
    .halt_o_t1(halt_ctrl_t1),
    .\resolved_branch_i.cf_type (\resolved_branch.cf_type ),
    .\resolved_branch_i.cf_type_t0 (\resolved_branch.cf_type_t0 ),
    .\resolved_branch_i.cf_type_t1 (\resolved_branch.cf_type_t1 ),
    .\resolved_branch_i.is_mispredict (\resolved_branch.is_mispredict ),
    .\resolved_branch_i.is_mispredict_t0 (\resolved_branch.is_mispredict_t0 ),
    .\resolved_branch_i.is_mispredict_t1 (\resolved_branch.is_mispredict_t1 ),
    .\resolved_branch_i.is_taken (\resolved_branch.is_taken ),
    .\resolved_branch_i.is_taken_t0 (\resolved_branch.is_taken_t0 ),
    .\resolved_branch_i.is_taken_t1 (\resolved_branch.is_taken_t1 ),
    .\resolved_branch_i.pc (\resolved_branch.pc ),
    .\resolved_branch_i.pc_t0 (\resolved_branch.pc_t0 ),
    .\resolved_branch_i.pc_t1 (\resolved_branch.pc_t1 ),
    .\resolved_branch_i.target_address (\resolved_branch.target_address ),
    .\resolved_branch_i.target_address_t0 (\resolved_branch.target_address_t0 ),
    .\resolved_branch_i.target_address_t1 (\resolved_branch.target_address_t1 ),
    .\resolved_branch_i.valid (\resolved_branch.valid ),
    .\resolved_branch_i.valid_t0 (\resolved_branch.valid_t0 ),
    .\resolved_branch_i.valid_t1 (\resolved_branch.valid_t1 ),
    .rst_ni(rst_ni),
    .set_debug_pc_i(set_debug_pc),
    .set_debug_pc_i_t0(set_debug_pc_t0),
    .set_debug_pc_i_t1(set_debug_pc_t1),
    .set_pc_commit_o(set_pc_ctrl_pcgen),
    .set_pc_commit_o_t0(set_pc_ctrl_pcgen_t0),
    .set_pc_commit_o_t1(set_pc_ctrl_pcgen_t1),
    .sfence_vma_i(sfence_vma_commit_controller),
    .sfence_vma_i_t0(sfence_vma_commit_controller_t0),
    .sfence_vma_i_t1(sfence_vma_commit_controller_t1)
  );
  \csr_regfile(AsidWidth=16,NrCommitPorts=32'b010,NrPMPEntries=32'b01000)  csr_regfile_i (
    .asid_o(asid_csr_ex),
    .asid_o_t0(asid_csr_ex_t0),
    .asid_o_t1(asid_csr_ex_t1),
    .boot_addr_i(64'h0000000000000000),
    .boot_addr_i_t0(64'h0000000000000000),
    .boot_addr_i_t1(64'h0000000000000000),
    .clk_i(clk_i),
    .commit_ack_i(commit_ack),
    .commit_ack_i_t0(commit_ack_t0),
    .commit_ack_i_t1(commit_ack_t1),
    .\commit_instr_i[0].bp.cf (\commit_instr_id_commit[0].bp.cf ),
    .\commit_instr_i[0].bp.cf_t0 (\commit_instr_id_commit[0].bp.cf_t0 ),
    .\commit_instr_i[0].bp.cf_t1 (\commit_instr_id_commit[0].bp.cf_t1 ),
    .\commit_instr_i[0].bp.predict_address (\commit_instr_id_commit[0].bp.predict_address ),
    .\commit_instr_i[0].bp.predict_address_t0 (\commit_instr_id_commit[0].bp.predict_address_t0 ),
    .\commit_instr_i[0].bp.predict_address_t1 (\commit_instr_id_commit[0].bp.predict_address_t1 ),
    .\commit_instr_i[0].ex.cause (\commit_instr_id_commit[0].ex.cause ),
    .\commit_instr_i[0].ex.cause_t0 (\commit_instr_id_commit[0].ex.cause_t0 ),
    .\commit_instr_i[0].ex.cause_t1 (\commit_instr_id_commit[0].ex.cause_t1 ),
    .\commit_instr_i[0].ex.tval (\commit_instr_id_commit[0].ex.tval ),
    .\commit_instr_i[0].ex.tval_t0 (\commit_instr_id_commit[0].ex.tval_t0 ),
    .\commit_instr_i[0].ex.tval_t1 (\commit_instr_id_commit[0].ex.tval_t1 ),
    .\commit_instr_i[0].ex.valid (\commit_instr_id_commit[0].ex.valid ),
    .\commit_instr_i[0].ex.valid_t0 (\commit_instr_id_commit[0].ex.valid_t0 ),
    .\commit_instr_i[0].ex.valid_t1 (\commit_instr_id_commit[0].ex.valid_t1 ),
    .\commit_instr_i[0].fu (\commit_instr_id_commit[0].fu ),
    .\commit_instr_i[0].fu_t0 (\commit_instr_id_commit[0].fu_t0 ),
    .\commit_instr_i[0].fu_t1 (\commit_instr_id_commit[0].fu_t1 ),
    .\commit_instr_i[0].is_compressed (\commit_instr_id_commit[0].is_compressed ),
    .\commit_instr_i[0].is_compressed_t0 (\commit_instr_id_commit[0].is_compressed_t0 ),
    .\commit_instr_i[0].is_compressed_t1 (\commit_instr_id_commit[0].is_compressed_t1 ),
    .\commit_instr_i[0].op (\commit_instr_id_commit[0].op ),
    .\commit_instr_i[0].op_t0 (\commit_instr_id_commit[0].op_t0 ),
    .\commit_instr_i[0].op_t1 (\commit_instr_id_commit[0].op_t1 ),
    .\commit_instr_i[0].pc (\commit_instr_id_commit[0].pc ),
    .\commit_instr_i[0].pc_t0 (\commit_instr_id_commit[0].pc_t0 ),
    .\commit_instr_i[0].pc_t1 (\commit_instr_id_commit[0].pc_t1 ),
    .\commit_instr_i[0].rd (\commit_instr_id_commit[0].rd ),
    .\commit_instr_i[0].rd_t0 (\commit_instr_id_commit[0].rd_t0 ),
    .\commit_instr_i[0].rd_t1 (\commit_instr_id_commit[0].rd_t1 ),
    .\commit_instr_i[0].result (\commit_instr_id_commit[0].result ),
    .\commit_instr_i[0].result_t0 (\commit_instr_id_commit[0].result_t0 ),
    .\commit_instr_i[0].result_t1 (\commit_instr_id_commit[0].result_t1 ),
    .\commit_instr_i[0].rs1 (\commit_instr_id_commit[0].rs1 ),
    .\commit_instr_i[0].rs1_t0 (\commit_instr_id_commit[0].rs1_t0 ),
    .\commit_instr_i[0].rs1_t1 (\commit_instr_id_commit[0].rs1_t1 ),
    .\commit_instr_i[0].rs2 (\commit_instr_id_commit[0].rs2 ),
    .\commit_instr_i[0].rs2_t0 (\commit_instr_id_commit[0].rs2_t0 ),
    .\commit_instr_i[0].rs2_t1 (\commit_instr_id_commit[0].rs2_t1 ),
    .\commit_instr_i[0].trans_id (\commit_instr_id_commit[0].trans_id ),
    .\commit_instr_i[0].trans_id_t0 (\commit_instr_id_commit[0].trans_id_t0 ),
    .\commit_instr_i[0].trans_id_t1 (\commit_instr_id_commit[0].trans_id_t1 ),
    .\commit_instr_i[0].use_imm (\commit_instr_id_commit[0].use_imm ),
    .\commit_instr_i[0].use_imm_t0 (\commit_instr_id_commit[0].use_imm_t0 ),
    .\commit_instr_i[0].use_imm_t1 (\commit_instr_id_commit[0].use_imm_t1 ),
    .\commit_instr_i[0].use_pc (\commit_instr_id_commit[0].use_pc ),
    .\commit_instr_i[0].use_pc_t0 (\commit_instr_id_commit[0].use_pc_t0 ),
    .\commit_instr_i[0].use_pc_t1 (\commit_instr_id_commit[0].use_pc_t1 ),
    .\commit_instr_i[0].use_zimm (\commit_instr_id_commit[0].use_zimm ),
    .\commit_instr_i[0].use_zimm_t0 (\commit_instr_id_commit[0].use_zimm_t0 ),
    .\commit_instr_i[0].use_zimm_t1 (\commit_instr_id_commit[0].use_zimm_t1 ),
    .\commit_instr_i[0].valid (\commit_instr_id_commit[0].valid ),
    .\commit_instr_i[0].valid_t0 (\commit_instr_id_commit[0].valid_t0 ),
    .\commit_instr_i[0].valid_t1 (\commit_instr_id_commit[0].valid_t1 ),
    .\commit_instr_i[1].bp.cf (\commit_instr_id_commit[1].bp.cf ),
    .\commit_instr_i[1].bp.cf_t0 (\commit_instr_id_commit[1].bp.cf_t0 ),
    .\commit_instr_i[1].bp.cf_t1 (\commit_instr_id_commit[1].bp.cf_t1 ),
    .\commit_instr_i[1].bp.predict_address (\commit_instr_id_commit[1].bp.predict_address ),
    .\commit_instr_i[1].bp.predict_address_t0 (\commit_instr_id_commit[1].bp.predict_address_t0 ),
    .\commit_instr_i[1].bp.predict_address_t1 (\commit_instr_id_commit[1].bp.predict_address_t1 ),
    .\commit_instr_i[1].ex.cause (\commit_instr_id_commit[1].ex.cause ),
    .\commit_instr_i[1].ex.cause_t0 (\commit_instr_id_commit[1].ex.cause_t0 ),
    .\commit_instr_i[1].ex.cause_t1 (\commit_instr_id_commit[1].ex.cause_t1 ),
    .\commit_instr_i[1].ex.tval (\commit_instr_id_commit[1].ex.tval ),
    .\commit_instr_i[1].ex.tval_t0 (\commit_instr_id_commit[1].ex.tval_t0 ),
    .\commit_instr_i[1].ex.tval_t1 (\commit_instr_id_commit[1].ex.tval_t1 ),
    .\commit_instr_i[1].ex.valid (\commit_instr_id_commit[1].ex.valid ),
    .\commit_instr_i[1].ex.valid_t0 (\commit_instr_id_commit[1].ex.valid_t0 ),
    .\commit_instr_i[1].ex.valid_t1 (\commit_instr_id_commit[1].ex.valid_t1 ),
    .\commit_instr_i[1].fu (\commit_instr_id_commit[1].fu ),
    .\commit_instr_i[1].fu_t0 (\commit_instr_id_commit[1].fu_t0 ),
    .\commit_instr_i[1].fu_t1 (\commit_instr_id_commit[1].fu_t1 ),
    .\commit_instr_i[1].is_compressed (\commit_instr_id_commit[1].is_compressed ),
    .\commit_instr_i[1].is_compressed_t0 (\commit_instr_id_commit[1].is_compressed_t0 ),
    .\commit_instr_i[1].is_compressed_t1 (\commit_instr_id_commit[1].is_compressed_t1 ),
    .\commit_instr_i[1].op (\commit_instr_id_commit[1].op ),
    .\commit_instr_i[1].op_t0 (\commit_instr_id_commit[1].op_t0 ),
    .\commit_instr_i[1].op_t1 (\commit_instr_id_commit[1].op_t1 ),
    .\commit_instr_i[1].pc (\commit_instr_id_commit[1].pc ),
    .\commit_instr_i[1].pc_t0 (\commit_instr_id_commit[1].pc_t0 ),
    .\commit_instr_i[1].pc_t1 (\commit_instr_id_commit[1].pc_t1 ),
    .\commit_instr_i[1].rd (\commit_instr_id_commit[1].rd ),
    .\commit_instr_i[1].rd_t0 (\commit_instr_id_commit[1].rd_t0 ),
    .\commit_instr_i[1].rd_t1 (\commit_instr_id_commit[1].rd_t1 ),
    .\commit_instr_i[1].result (\commit_instr_id_commit[1].result ),
    .\commit_instr_i[1].result_t0 (\commit_instr_id_commit[1].result_t0 ),
    .\commit_instr_i[1].result_t1 (\commit_instr_id_commit[1].result_t1 ),
    .\commit_instr_i[1].rs1 (\commit_instr_id_commit[1].rs1 ),
    .\commit_instr_i[1].rs1_t0 (\commit_instr_id_commit[1].rs1_t0 ),
    .\commit_instr_i[1].rs1_t1 (\commit_instr_id_commit[1].rs1_t1 ),
    .\commit_instr_i[1].rs2 (\commit_instr_id_commit[1].rs2 ),
    .\commit_instr_i[1].rs2_t0 (\commit_instr_id_commit[1].rs2_t0 ),
    .\commit_instr_i[1].rs2_t1 (\commit_instr_id_commit[1].rs2_t1 ),
    .\commit_instr_i[1].trans_id (\commit_instr_id_commit[1].trans_id ),
    .\commit_instr_i[1].trans_id_t0 (\commit_instr_id_commit[1].trans_id_t0 ),
    .\commit_instr_i[1].trans_id_t1 (\commit_instr_id_commit[1].trans_id_t1 ),
    .\commit_instr_i[1].use_imm (\commit_instr_id_commit[1].use_imm ),
    .\commit_instr_i[1].use_imm_t0 (\commit_instr_id_commit[1].use_imm_t0 ),
    .\commit_instr_i[1].use_imm_t1 (\commit_instr_id_commit[1].use_imm_t1 ),
    .\commit_instr_i[1].use_pc (\commit_instr_id_commit[1].use_pc ),
    .\commit_instr_i[1].use_pc_t0 (\commit_instr_id_commit[1].use_pc_t0 ),
    .\commit_instr_i[1].use_pc_t1 (\commit_instr_id_commit[1].use_pc_t1 ),
    .\commit_instr_i[1].use_zimm (\commit_instr_id_commit[1].use_zimm ),
    .\commit_instr_i[1].use_zimm_t0 (\commit_instr_id_commit[1].use_zimm_t0 ),
    .\commit_instr_i[1].use_zimm_t1 (\commit_instr_id_commit[1].use_zimm_t1 ),
    .\commit_instr_i[1].valid (\commit_instr_id_commit[1].valid ),
    .\commit_instr_i[1].valid_t0 (\commit_instr_id_commit[1].valid_t0 ),
    .\commit_instr_i[1].valid_t1 (\commit_instr_id_commit[1].valid_t1 ),
    .csr_addr_i(csr_addr_ex_csr),
    .csr_addr_i_t0(csr_addr_ex_csr_t0),
    .csr_addr_i_t1(csr_addr_ex_csr_t1),
    .\csr_exception_o.cause (\csr_exception_csr_commit.cause ),
    .\csr_exception_o.cause_t0 (\csr_exception_csr_commit.cause_t0 ),
    .\csr_exception_o.cause_t1 (\csr_exception_csr_commit.cause_t1 ),
    .\csr_exception_o.tval (\csr_exception_csr_commit.tval ),
    .\csr_exception_o.tval_t0 (\csr_exception_csr_commit.tval_t0 ),
    .\csr_exception_o.tval_t1 (\csr_exception_csr_commit.tval_t1 ),
    .\csr_exception_o.valid (\csr_exception_csr_commit.valid ),
    .\csr_exception_o.valid_t0 (\csr_exception_csr_commit.valid_t0 ),
    .\csr_exception_o.valid_t1 (\csr_exception_csr_commit.valid_t1 ),
    .csr_op_i(csr_op_commit_csr),
    .csr_op_i_t0(csr_op_commit_csr_t0),
    .csr_op_i_t1(csr_op_commit_csr_t1),
    .csr_rdata_o(csr_rdata_csr_commit),
    .csr_rdata_o_t0(csr_rdata_csr_commit_t0),
    .csr_rdata_o_t1(csr_rdata_csr_commit_t1),
    .csr_wdata_i(csr_wdata_commit_csr),
    .csr_wdata_i_t0(csr_wdata_commit_csr_t0),
    .csr_wdata_i_t1(csr_wdata_commit_csr_t1),
    .csr_write_fflags_i(csr_write_fflags_commit_cs),
    .csr_write_fflags_i_t0(csr_write_fflags_commit_cs_t0),
    .csr_write_fflags_i_t1(csr_write_fflags_commit_cs_t1),
    .dcache_en_o(dcache_en_csr_nbdcache),
    .dcache_en_o_t0(dcache_en_csr_nbdcache_t0),
    .dcache_en_o_t1(dcache_en_csr_nbdcache_t1),
    .debug_mode_o(debug_mode),
    .debug_mode_o_t0(debug_mode_t0),
    .debug_mode_o_t1(debug_mode_t1),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .debug_req_i_t1(debug_req_i_t1),
    .dirty_fp_state_i(dirty_fp_state),
    .dirty_fp_state_i_t0(dirty_fp_state_t0),
    .dirty_fp_state_i_t1(dirty_fp_state_t1),
    .en_ld_st_translation_o(en_ld_st_translation_csr_ex),
    .en_ld_st_translation_o_t0(en_ld_st_translation_csr_ex_t0),
    .en_ld_st_translation_o_t1(en_ld_st_translation_csr_ex_t1),
    .en_translation_o(enable_translation_csr_ex),
    .en_translation_o_t0(enable_translation_csr_ex_t0),
    .en_translation_o_t1(enable_translation_csr_ex_t1),
    .epc_o(epc_commit_pcgen),
    .epc_o_t0(epc_commit_pcgen_t0),
    .epc_o_t1(epc_commit_pcgen_t1),
    .eret_o(eret),
    .eret_o_t0(eret_t0),
    .eret_o_t1(eret_t1),
    .\ex_i.cause (\ex_commit.cause ),
    .\ex_i.cause_t0 (\ex_commit.cause_t0 ),
    .\ex_i.cause_t1 (\ex_commit.cause_t1 ),
    .\ex_i.tval (\ex_commit.tval ),
    .\ex_i.tval_t0 (\ex_commit.tval_t0 ),
    .\ex_i.tval_t1 (\ex_commit.tval_t1 ),
    .\ex_i.valid (\ex_commit.valid ),
    .\ex_i.valid_t0 (\ex_commit.valid_t0 ),
    .\ex_i.valid_t1 (\ex_commit.valid_t1 ),
    .fflags_o(fflags_csr_commit),
    .fflags_o_t0(fflags_csr_commit_t0),
    .fflags_o_t1(fflags_csr_commit_t1),
    .flush_o(flush_csr_ctrl),
    .flush_o_t0(flush_csr_ctrl_t0),
    .flush_o_t1(flush_csr_ctrl_t1),
    .fprec_o(fprec_csr_ex),
    .fprec_o_t0(fprec_csr_ex_t0),
    .fprec_o_t1(fprec_csr_ex_t1),
    .frm_o(frm_csr_id_issue_ex),
    .frm_o_t0(frm_csr_id_issue_ex_t0),
    .frm_o_t1(frm_csr_id_issue_ex_t1),
    .fs_o(fs),
    .fs_o_t0(fs_t0),
    .fs_o_t1(fs_t1),
    .halt_csr_o(halt_csr_ctrl),
    .halt_csr_o_t0(halt_csr_ctrl_t0),
    .halt_csr_o_t1(halt_csr_ctrl_t1),
    .hart_id_i(64'h0000000000000000),
    .hart_id_i_t0(64'h0000000000000000),
    .hart_id_i_t1(64'h0000000000000000),
    .icache_en_o(icache_en_csr),
    .icache_en_o_t0(icache_en_csr_t0),
    .icache_en_o_t1(icache_en_csr_t1),
    .ipi_i(ipi_i),
    .ipi_i_t0(ipi_i_t0),
    .ipi_i_t1(ipi_i_t1),
    .\irq_ctrl_o.global_enable (\irq_ctrl_csr_id.global_enable ),
    .\irq_ctrl_o.global_enable_t0 (\irq_ctrl_csr_id.global_enable_t0 ),
    .\irq_ctrl_o.global_enable_t1 (\irq_ctrl_csr_id.global_enable_t1 ),
    .\irq_ctrl_o.mideleg (\irq_ctrl_csr_id.mideleg ),
    .\irq_ctrl_o.mideleg_t0 (\irq_ctrl_csr_id.mideleg_t0 ),
    .\irq_ctrl_o.mideleg_t1 (\irq_ctrl_csr_id.mideleg_t1 ),
    .\irq_ctrl_o.mie (\irq_ctrl_csr_id.mie ),
    .\irq_ctrl_o.mie_t0 (\irq_ctrl_csr_id.mie_t0 ),
    .\irq_ctrl_o.mie_t1 (\irq_ctrl_csr_id.mie_t1 ),
    .\irq_ctrl_o.mip (\irq_ctrl_csr_id.mip ),
    .\irq_ctrl_o.mip_t0 (\irq_ctrl_csr_id.mip_t0 ),
    .\irq_ctrl_o.mip_t1 (\irq_ctrl_csr_id.mip_t1 ),
    .\irq_ctrl_o.sie (\irq_ctrl_csr_id.sie ),
    .\irq_ctrl_o.sie_t0 (\irq_ctrl_csr_id.sie_t0 ),
    .\irq_ctrl_o.sie_t1 (\irq_ctrl_csr_id.sie_t1 ),
    .irq_i(2'h0),
    .irq_i_t0(2'h0),
    .irq_i_t1(2'h0),
    .ld_st_priv_lvl_o(ld_st_priv_lvl_csr_ex),
    .ld_st_priv_lvl_o_t0(ld_st_priv_lvl_csr_ex_t0),
    .ld_st_priv_lvl_o_t1(ld_st_priv_lvl_csr_ex_t1),
    .mxr_o(mxr_csr_ex),
    .mxr_o_t0(mxr_csr_ex_t0),
    .mxr_o_t1(mxr_csr_ex_t1),
    .pc_i(pc_commit),
    .pc_i_t0(pc_commit_t0),
    .pc_i_t1(pc_commit_t1),
    .priv_lvl_o(priv_lvl),
    .priv_lvl_o_t0(priv_lvl_t0),
    .priv_lvl_o_t1(priv_lvl_t1),
    .rst_ni(rst_ni),
    .satp_ppn_o(satp_ppn_csr_ex),
    .satp_ppn_o_t0(satp_ppn_csr_ex_t0),
    .satp_ppn_o_t1(satp_ppn_csr_ex_t1),
    .set_debug_pc_o(set_debug_pc),
    .set_debug_pc_o_t0(set_debug_pc_t0),
    .set_debug_pc_o_t1(set_debug_pc_t1),
    .single_step_o(single_step_csr_commit),
    .single_step_o_t0(single_step_csr_commit_t0),
    .single_step_o_t1(single_step_csr_commit_t1),
    .sum_o(sum_csr_ex),
    .sum_o_t0(sum_csr_ex_t0),
    .sum_o_t1(sum_csr_ex_t1),
    .time_irq_i(time_irq_i),
    .time_irq_i_t0(time_irq_i_t0),
    .time_irq_i_t1(time_irq_i_t1),
    .trap_vector_base_o(trap_vector_base_commit_pcgen),
    .trap_vector_base_o_t0(trap_vector_base_commit_pcgen_t0),
    .trap_vector_base_o_t1(trap_vector_base_commit_pcgen_t1),
    .tsr_o(tsr_csr_id),
    .tsr_o_t0(tsr_csr_id_t0),
    .tsr_o_t1(tsr_csr_id_t1),
    .tvm_o(tvm_csr_id),
    .tvm_o_t0(tvm_csr_id_t0),
    .tvm_o_t1(tvm_csr_id_t1),
    .tw_o(tw_csr_id),
    .tw_o_t0(tw_csr_id_t0),
    .tw_o_t1(tw_csr_id_t1)
  );
  \ex_stage(ASID_WIDTH=32'b010000,ArianeCfg='{2,32,128,32'b010,1024'b0,1024'b0,32'b011,1024'b01000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000,1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000,32'b01,1024'b010000000000000000000000000000000,1024'b01000000000000000000000000000000,1'b1,1'b0,64'b0,32'b01000})  ex_stage_i (
    .alu_valid_i(alu_valid_id_ex),
    .alu_valid_i_t0(alu_valid_id_ex_t0),
    .alu_valid_i_t1(alu_valid_id_ex_t1),
    .amo_valid_commit_i(amo_valid_commit),
    .amo_valid_commit_i_t0(amo_valid_commit_t0),
    .amo_valid_commit_i_t1(amo_valid_commit_t1),
    .asid_i(asid_csr_ex),
    .asid_i_t0(asid_csr_ex_t0),
    .asid_i_t1(asid_csr_ex_t1),
    .\branch_predict_i.cf (\branch_predict_id_ex.cf ),
    .\branch_predict_i.cf_t0 (\branch_predict_id_ex.cf_t0 ),
    .\branch_predict_i.cf_t1 (\branch_predict_id_ex.cf_t1 ),
    .\branch_predict_i.predict_address (\branch_predict_id_ex.predict_address ),
    .\branch_predict_i.predict_address_t0 (\branch_predict_id_ex.predict_address_t0 ),
    .\branch_predict_i.predict_address_t1 (\branch_predict_id_ex.predict_address_t1 ),
    .branch_valid_i(branch_valid_id_ex),
    .branch_valid_i_t0(branch_valid_id_ex_t0),
    .branch_valid_i_t1(branch_valid_id_ex_t1),
    .clk_i(clk_i),
    .commit_tran_id_i(lsu_commit_trans_id),
    .commit_tran_id_i_t0(lsu_commit_trans_id_t0),
    .commit_tran_id_i_t1(lsu_commit_trans_id_t1),
    .csr_addr_o(csr_addr_ex_csr),
    .csr_addr_o_t0(csr_addr_ex_csr_t0),
    .csr_addr_o_t1(csr_addr_ex_csr_t1),
    .csr_commit_i(csr_commit_commit_ex),
    .csr_commit_i_t0(csr_commit_commit_ex_t0),
    .csr_commit_i_t1(csr_commit_commit_ex_t1),
    .csr_valid_i(csr_valid_id_ex),
    .csr_valid_i_t0(csr_valid_id_ex_t0),
    .csr_valid_i_t1(csr_valid_id_ex_t1),
    .debug_mode_i(debug_mode),
    .debug_mode_i_t0(debug_mode_t0),
    .debug_mode_i_t1(debug_mode_t1),
    .en_ld_st_translation_i(en_ld_st_translation_csr_ex),
    .en_ld_st_translation_i_t0(en_ld_st_translation_csr_ex_t0),
    .en_ld_st_translation_i_t1(en_ld_st_translation_csr_ex_t1),
    .enable_translation_i(enable_translation_csr_ex),
    .enable_translation_i_t0(enable_translation_csr_ex_t0),
    .enable_translation_i_t1(enable_translation_csr_ex_t1),
    .\flu_exception_o.cause (\flu_exception_ex_id.cause ),
    .\flu_exception_o.cause_t0 (\flu_exception_ex_id.cause_t0 ),
    .\flu_exception_o.cause_t1 (\flu_exception_ex_id.cause_t1 ),
    .\flu_exception_o.tval (\flu_exception_ex_id.tval ),
    .\flu_exception_o.tval_t0 (\flu_exception_ex_id.tval_t0 ),
    .\flu_exception_o.tval_t1 (\flu_exception_ex_id.tval_t1 ),
    .\flu_exception_o.valid (\flu_exception_ex_id.valid ),
    .\flu_exception_o.valid_t0 (\flu_exception_ex_id.valid_t0 ),
    .\flu_exception_o.valid_t1 (\flu_exception_ex_id.valid_t1 ),
    .flu_ready_o(flu_ready_ex_id),
    .flu_ready_o_t0(flu_ready_ex_id_t0),
    .flu_ready_o_t1(flu_ready_ex_id_t1),
    .flu_result_o(flu_result_ex_id),
    .flu_result_o_t0(flu_result_ex_id_t0),
    .flu_result_o_t1(flu_result_ex_id_t1),
    .flu_trans_id_o(flu_trans_id_ex_id),
    .flu_trans_id_o_t0(flu_trans_id_ex_id_t0),
    .flu_trans_id_o_t1(flu_trans_id_ex_id_t1),
    .flu_valid_o(flu_valid_ex_id),
    .flu_valid_o_t0(flu_valid_ex_id_t0),
    .flu_valid_o_t1(flu_valid_ex_id_t1),
    .flush_i(flush_ctrl_ex),
    .flush_i_t0(flush_ctrl_ex_t0),
    .flush_i_t1(flush_ctrl_ex_t1),
    .flush_tlb_i(flush_tlb_ctrl_ex),
    .flush_tlb_i_t0(flush_tlb_ctrl_ex_t0),
    .flush_tlb_i_t1(flush_tlb_ctrl_ex_t1),
    .\fpu_exception_o.cause (\fpu_exception_ex_id.cause ),
    .\fpu_exception_o.cause_t0 (\fpu_exception_ex_id.cause_t0 ),
    .\fpu_exception_o.cause_t1 (\fpu_exception_ex_id.cause_t1 ),
    .\fpu_exception_o.tval (\fpu_exception_ex_id.tval ),
    .\fpu_exception_o.tval_t0 (\fpu_exception_ex_id.tval_t0 ),
    .\fpu_exception_o.tval_t1 (\fpu_exception_ex_id.tval_t1 ),
    .\fpu_exception_o.valid (\fpu_exception_ex_id.valid ),
    .\fpu_exception_o.valid_t0 (\fpu_exception_ex_id.valid_t0 ),
    .\fpu_exception_o.valid_t1 (\fpu_exception_ex_id.valid_t1 ),
    .fpu_fmt_i(fpu_fmt_id_ex),
    .fpu_fmt_i_t0(fpu_fmt_id_ex_t0),
    .fpu_fmt_i_t1(fpu_fmt_id_ex_t1),
    .fpu_frm_i(frm_csr_id_issue_ex),
    .fpu_frm_i_t0(frm_csr_id_issue_ex_t0),
    .fpu_frm_i_t1(frm_csr_id_issue_ex_t1),
    .fpu_prec_i(fprec_csr_ex),
    .fpu_prec_i_t0(fprec_csr_ex_t0),
    .fpu_prec_i_t1(fprec_csr_ex_t1),
    .fpu_ready_o(fpu_ready_ex_id),
    .fpu_ready_o_t0(fpu_ready_ex_id_t0),
    .fpu_ready_o_t1(fpu_ready_ex_id_t1),
    .fpu_result_o(fpu_result_ex_id),
    .fpu_result_o_t0(fpu_result_ex_id_t0),
    .fpu_result_o_t1(fpu_result_ex_id_t1),
    .fpu_rm_i(fpu_rm_id_ex),
    .fpu_rm_i_t0(fpu_rm_id_ex_t0),
    .fpu_rm_i_t1(fpu_rm_id_ex_t1),
    .fpu_trans_id_o(fpu_trans_id_ex_id),
    .fpu_trans_id_o_t0(fpu_trans_id_ex_id_t0),
    .fpu_trans_id_o_t1(fpu_trans_id_ex_id_t1),
    .fpu_valid_i(fpu_valid_id_ex),
    .fpu_valid_i_t0(fpu_valid_id_ex_t0),
    .fpu_valid_i_t1(fpu_valid_id_ex_t1),
    .fpu_valid_o(fpu_valid_ex_id),
    .fpu_valid_o_t0(fpu_valid_ex_id_t0),
    .fpu_valid_o_t1(fpu_valid_ex_id_t1),
    .\fu_data_i.fu (\fu_data_id_ex.fu ),
    .\fu_data_i.fu_t0 (\fu_data_id_ex.fu_t0 ),
    .\fu_data_i.fu_t1 (\fu_data_id_ex.fu_t1 ),
    .\fu_data_i.imm (\fu_data_id_ex.imm ),
    .\fu_data_i.imm_t0 (\fu_data_id_ex.imm_t0 ),
    .\fu_data_i.imm_t1 (\fu_data_id_ex.imm_t1 ),
    .\fu_data_i.operand_a (\fu_data_id_ex.operand_a ),
    .\fu_data_i.operand_a_t0 (\fu_data_id_ex.operand_a_t0 ),
    .\fu_data_i.operand_a_t1 (\fu_data_id_ex.operand_a_t1 ),
    .\fu_data_i.operand_b (\fu_data_id_ex.operand_b ),
    .\fu_data_i.operand_b_t0 (\fu_data_id_ex.operand_b_t0 ),
    .\fu_data_i.operand_b_t1 (\fu_data_id_ex.operand_b_t1 ),
    .\fu_data_i.operator (\fu_data_id_ex.operator ),
    .\fu_data_i.operator_t0 (\fu_data_id_ex.operator_t0 ),
    .\fu_data_i.operator_t1 (\fu_data_id_ex.operator_t1 ),
    .\fu_data_i.trans_id (\fu_data_id_ex.trans_id ),
    .\fu_data_i.trans_id_t0 (\fu_data_id_ex.trans_id_t0 ),
    .\fu_data_i.trans_id_t1 (\fu_data_id_ex.trans_id_t1 ),
    .is_compressed_instr_i(is_compressed_instr_id_ex),
    .is_compressed_instr_i_t0(is_compressed_instr_id_ex_t0),
    .is_compressed_instr_i_t1(is_compressed_instr_id_ex_t1),
    .ld_st_priv_lvl_i(ld_st_priv_lvl_csr_ex),
    .ld_st_priv_lvl_i_t0(ld_st_priv_lvl_csr_ex_t0),
    .ld_st_priv_lvl_i_t1(ld_st_priv_lvl_csr_ex_t1),
    .\load_exception_o.cause (\load_exception_ex_id.cause ),
    .\load_exception_o.cause_t0 (\load_exception_ex_id.cause_t0 ),
    .\load_exception_o.cause_t1 (\load_exception_ex_id.cause_t1 ),
    .\load_exception_o.tval (\load_exception_ex_id.tval ),
    .\load_exception_o.tval_t0 (\load_exception_ex_id.tval_t0 ),
    .\load_exception_o.tval_t1 (\load_exception_ex_id.tval_t1 ),
    .\load_exception_o.valid (\load_exception_ex_id.valid ),
    .\load_exception_o.valid_t0 (\load_exception_ex_id.valid_t0 ),
    .\load_exception_o.valid_t1 (\load_exception_ex_id.valid_t1 ),
    .load_result_o(load_result_ex_id),
    .load_result_o_t0(load_result_ex_id_t0),
    .load_result_o_t1(load_result_ex_id_t1),
    .load_trans_id_o(load_trans_id_ex_id),
    .load_trans_id_o_t0(load_trans_id_ex_id_t0),
    .load_trans_id_o_t1(load_trans_id_ex_id_t1),
    .load_valid_o(load_valid_ex_id),
    .load_valid_o_t0(load_valid_ex_id_t0),
    .load_valid_o_t1(load_valid_ex_id_t1),
    .lsu_commit_i(lsu_commit_commit_ex),
    .lsu_commit_i_t0(lsu_commit_commit_ex_t0),
    .lsu_commit_i_t1(lsu_commit_commit_ex_t1),
    .lsu_commit_ready_o(lsu_commit_ready_ex_commit),
    .lsu_commit_ready_o_t0(lsu_commit_ready_ex_commit_t0),
    .lsu_commit_ready_o_t1(lsu_commit_ready_ex_commit_t1),
    .lsu_ready_o(lsu_ready_ex_id),
    .lsu_ready_o_t0(lsu_ready_ex_id_t0),
    .lsu_ready_o_t1(lsu_ready_ex_id_t1),
    .lsu_valid_i(lsu_valid_id_ex),
    .lsu_valid_i_t0(lsu_valid_id_ex_t0),
    .lsu_valid_i_t1(lsu_valid_id_ex_t1),
    .mult_valid_i(mult_valid_id_ex),
    .mult_valid_i_t0(mult_valid_id_ex_t0),
    .mult_valid_i_t1(mult_valid_id_ex_t1),
    .mxr_i(mxr_csr_ex),
    .mxr_i_t0(mxr_csr_ex_t0),
    .mxr_i_t1(mxr_csr_ex_t1),
    .no_st_pending_o(no_st_pending_ex),
    .no_st_pending_o_t0(no_st_pending_ex_t0),
    .no_st_pending_o_t1(no_st_pending_ex_t1),
    .pc_i(pc_id_ex),
    .pc_i_t0(pc_id_ex_t0),
    .pc_i_t1(pc_id_ex_t1),
    .priv_lvl_i(priv_lvl),
    .priv_lvl_i_t0(priv_lvl_t0),
    .priv_lvl_i_t1(priv_lvl_t1),
    .resolve_branch_o(resolve_branch_ex_id),
    .resolve_branch_o_t0(resolve_branch_ex_id_t0),
    .resolve_branch_o_t1(resolve_branch_ex_id_t1),
    .\resolved_branch_o.cf_type (\resolved_branch.cf_type ),
    .\resolved_branch_o.cf_type_t0 (\resolved_branch.cf_type_t0 ),
    .\resolved_branch_o.cf_type_t1 (\resolved_branch.cf_type_t1 ),
    .\resolved_branch_o.is_mispredict (\resolved_branch.is_mispredict ),
    .\resolved_branch_o.is_mispredict_t0 (\resolved_branch.is_mispredict_t0 ),
    .\resolved_branch_o.is_mispredict_t1 (\resolved_branch.is_mispredict_t1 ),
    .\resolved_branch_o.is_taken (\resolved_branch.is_taken ),
    .\resolved_branch_o.is_taken_t0 (\resolved_branch.is_taken_t0 ),
    .\resolved_branch_o.is_taken_t1 (\resolved_branch.is_taken_t1 ),
    .\resolved_branch_o.pc (\resolved_branch.pc ),
    .\resolved_branch_o.pc_t0 (\resolved_branch.pc_t0 ),
    .\resolved_branch_o.pc_t1 (\resolved_branch.pc_t1 ),
    .\resolved_branch_o.target_address (\resolved_branch.target_address ),
    .\resolved_branch_o.target_address_t0 (\resolved_branch.target_address_t0 ),
    .\resolved_branch_o.target_address_t1 (\resolved_branch.target_address_t1 ),
    .\resolved_branch_o.valid (\resolved_branch.valid ),
    .\resolved_branch_o.valid_t0 (\resolved_branch.valid_t0 ),
    .\resolved_branch_o.valid_t1 (\resolved_branch.valid_t1 ),
    .rs1_forwarding_i(rs1_forwarding_id_ex),
    .rs1_forwarding_i_t0(rs1_forwarding_id_ex_t0),
    .rs1_forwarding_i_t1(rs1_forwarding_id_ex_t1),
    .rs2_forwarding_i(rs2_forwarding_id_ex),
    .rs2_forwarding_i_t0(rs2_forwarding_id_ex_t0),
    .rs2_forwarding_i_t1(rs2_forwarding_id_ex_t1),
    .rst_ni(rst_ni),
    .satp_ppn_i(satp_ppn_csr_ex),
    .satp_ppn_i_t0(satp_ppn_csr_ex_t0),
    .satp_ppn_i_t1(satp_ppn_csr_ex_t1),
    .\store_exception_o.cause (\store_exception_ex_id.cause ),
    .\store_exception_o.cause_t0 (\store_exception_ex_id.cause_t0 ),
    .\store_exception_o.cause_t1 (\store_exception_ex_id.cause_t1 ),
    .\store_exception_o.tval (\store_exception_ex_id.tval ),
    .\store_exception_o.tval_t0 (\store_exception_ex_id.tval_t0 ),
    .\store_exception_o.tval_t1 (\store_exception_ex_id.tval_t1 ),
    .\store_exception_o.valid (\store_exception_ex_id.valid ),
    .\store_exception_o.valid_t0 (\store_exception_ex_id.valid_t0 ),
    .\store_exception_o.valid_t1 (\store_exception_ex_id.valid_t1 ),
    .store_result_o(store_result_ex_id),
    .store_result_o_t0(store_result_ex_id_t0),
    .store_result_o_t1(store_result_ex_id_t1),
    .store_trans_id_o(store_trans_id_ex_id),
    .store_trans_id_o_t0(store_trans_id_ex_id_t0),
    .store_trans_id_o_t1(store_trans_id_ex_id_t1),
    .store_valid_o(store_valid_ex_id),
    .store_valid_o_t0(store_valid_ex_id_t0),
    .store_valid_o_t1(store_valid_ex_id_t1),
    .sum_i(sum_csr_ex),
    .sum_i_t0(sum_csr_ex_t0),
    .sum_i_t1(sum_csr_ex_t1)
  );
  //\frontend(ArianeCfg='{2,32,128,32'b010,1024'b0,1024'b0,32'b011,1024'b01000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000,1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000,32'b01,1024'b010000000000000000000000000000000,1024'b01000000000000000000000000000000,1'b1,1'b0,64'b0,32'b01000})  i_frontend (
  //  .boot_addr_i(64'h0000000000000000),
  //  .boot_addr_i_t0(64'h0000000000000000),
  //  .boot_addr_i_t1(64'h0000000000000000),
  //  .clk_i(clk_i),
  //  .debug_mode_i(debug_mode),
  //  .debug_mode_i_t0(debug_mode_t0),
  //  .debug_mode_i_t1(debug_mode_t1),
  //  .epc_i(epc_commit_pcgen),
  //  .epc_i_t0(epc_commit_pcgen_t0),
  //  .epc_i_t1(epc_commit_pcgen_t1),
  //  .eret_i(eret),
  //  .eret_i_t0(eret_t0),
  //  .eret_i_t1(eret_t1),
  //  .ex_valid_i(\ex_commit.valid ),
  //  .ex_valid_i_t0(\ex_commit.valid_t0 ),
  //  .ex_valid_i_t1(\ex_commit.valid_t1 ),
  //  .\fetch_entry_o.address (\fetch_entry_if_id.address ),
  //  .\fetch_entry_o.address_t0 (\fetch_entry_if_id.address_t0 ),
  //  .\fetch_entry_o.address_t1 (\fetch_entry_if_id.address_t1 ),
  //  .\fetch_entry_o.branch_predict.cf (\fetch_entry_if_id.branch_predict.cf ),
  //  .\fetch_entry_o.branch_predict.cf_t0 (\fetch_entry_if_id.branch_predict.cf_t0 ),
  //  .\fetch_entry_o.branch_predict.cf_t1 (\fetch_entry_if_id.branch_predict.cf_t1 ),
  //  .\fetch_entry_o.branch_predict.predict_address (\fetch_entry_if_id.branch_predict.predict_address ),
  //  .\fetch_entry_o.branch_predict.predict_address_t0 (\fetch_entry_if_id.branch_predict.predict_address_t0 ),
  //  .\fetch_entry_o.branch_predict.predict_address_t1 (\fetch_entry_if_id.branch_predict.predict_address_t1 ),
  //  .\fetch_entry_o.ex.cause (\fetch_entry_if_id.ex.cause ),
  //  .\fetch_entry_o.ex.cause_t0 (\fetch_entry_if_id.ex.cause_t0 ),
  //  .\fetch_entry_o.ex.cause_t1 (\fetch_entry_if_id.ex.cause_t1 ),
  //  .\fetch_entry_o.ex.tval (\fetch_entry_if_id.ex.tval ),
  //  .\fetch_entry_o.ex.tval_t0 (\fetch_entry_if_id.ex.tval_t0 ),
  //  .\fetch_entry_o.ex.tval_t1 (\fetch_entry_if_id.ex.tval_t1 ),
  //  .\fetch_entry_o.ex.valid (\fetch_entry_if_id.ex.valid ),
  //  .\fetch_entry_o.ex.valid_t0 (\fetch_entry_if_id.ex.valid_t0 ),
  //  .\fetch_entry_o.ex.valid_t1 (\fetch_entry_if_id.ex.valid_t1 ),
  //  .\fetch_entry_o.instruction (\fetch_entry_if_id.instruction ),
  //  .\fetch_entry_o.instruction_t0 (\fetch_entry_if_id.instruction_t0 ),
  //  .\fetch_entry_o.instruction_t1 (\fetch_entry_if_id.instruction_t1 ),
  //  .fetch_entry_ready_i(fetch_ready_id_if),
  //  .fetch_entry_ready_i_t0(fetch_ready_id_if_t0),
  //  .fetch_entry_ready_i_t1(fetch_ready_id_if_t1),
  //  .fetch_entry_valid_o(fetch_valid_if_id),
  //  .fetch_entry_valid_o_t0(fetch_valid_if_id_t0),
  //  .fetch_entry_valid_o_t1(fetch_valid_if_id_t1),
  //  .flush_bp_i(1'h0),
  //  .flush_bp_i_t0(1'h0),
  //  .flush_bp_i_t1(1'h0),
  //  .flush_i(flush_ctrl_if),
  //  .flush_i_t0(flush_ctrl_if_t0),
  //  .flush_i_t1(flush_ctrl_if_t1),
  //  .\icache_dreq_i.data (\tmp_icache_dreq_cache_if.data ),
  //  .\icache_dreq_i.data_t0 (\tmp_icache_dreq_cache_if.data_t0 ),
  //  .\icache_dreq_i.data_t1 (\tmp_icache_dreq_cache_if.data_t1 ),
  //  .\icache_dreq_i.ex.cause (\tmp_icache_dreq_cache_if.ex.cause ),
  //  .\icache_dreq_i.ex.cause_t0 (\tmp_icache_dreq_cache_if.ex.cause_t0 ),
  //  .\icache_dreq_i.ex.cause_t1 (\tmp_icache_dreq_cache_if.ex.cause_t1 ),
  //  .\icache_dreq_i.ex.tval (\tmp_icache_dreq_cache_if.ex.tval ),
  //  .\icache_dreq_i.ex.tval_t0 (\tmp_icache_dreq_cache_if.ex.tval_t0 ),
  //  .\icache_dreq_i.ex.tval_t1 (\tmp_icache_dreq_cache_if.ex.tval_t1 ),
  //  .\icache_dreq_i.ex.valid (\tmp_icache_dreq_cache_if.ex.valid ),
  //  .\icache_dreq_i.ex.valid_t0 (\tmp_icache_dreq_cache_if.ex.valid_t0 ),
  //  .\icache_dreq_i.ex.valid_t1 (\tmp_icache_dreq_cache_if.ex.valid_t1 ),
  //  .\icache_dreq_i.ready (\tmp_icache_dreq_cache_if.ready ),
  //  .\icache_dreq_i.ready_t0 (\tmp_icache_dreq_cache_if.ready_t0 ),
  //  .\icache_dreq_i.ready_t1 (\tmp_icache_dreq_cache_if.ready_t1 ),
  //  .\icache_dreq_i.vaddr (\tmp_icache_dreq_cache_if.vaddr ),
  //  .\icache_dreq_i.vaddr_t0 (\tmp_icache_dreq_cache_if.vaddr_t0 ),
  //  .\icache_dreq_i.vaddr_t1 (\tmp_icache_dreq_cache_if.vaddr_t1 ),
  //  .\icache_dreq_i.valid (\tmp_icache_dreq_cache_if.valid ),
  //  .\icache_dreq_i.valid_t0 (\tmp_icache_dreq_cache_if.valid_t0 ),
  //  .\icache_dreq_i.valid_t1 (\tmp_icache_dreq_cache_if.valid_t1 ),
  //  .\icache_dreq_o.kill_s1 (\tmp_icache_dreq_if_cache.kill_s1 ),
  //  .\icache_dreq_o.kill_s1_t0 (\tmp_icache_dreq_if_cache.kill_s1_t0 ),
  //  .\icache_dreq_o.kill_s1_t1 (\tmp_icache_dreq_if_cache.kill_s1_t1 ),
  //  .\icache_dreq_o.kill_s2 (\tmp_icache_dreq_if_cache.kill_s2 ),
  //  .\icache_dreq_o.kill_s2_t0 (\tmp_icache_dreq_if_cache.kill_s2_t0 ),
  //  .\icache_dreq_o.kill_s2_t1 (\tmp_icache_dreq_if_cache.kill_s2_t1 ),
  //  .\icache_dreq_o.req (\tmp_icache_dreq_if_cache.req ),
  //  .\icache_dreq_o.req_t0 (\tmp_icache_dreq_if_cache.req_t0 ),
  //  .\icache_dreq_o.req_t1 (\tmp_icache_dreq_if_cache.req_t1 ),
  //  .\icache_dreq_o.spec (\tmp_icache_dreq_if_cache.spec ),
  //  .\icache_dreq_o.spec_t0 (\tmp_icache_dreq_if_cache.spec_t0 ),
  //  .\icache_dreq_o.spec_t1 (\tmp_icache_dreq_if_cache.spec_t1 ),
  //  .\icache_dreq_o.vaddr (\tmp_icache_dreq_if_cache.vaddr ),
  //  .\icache_dreq_o.vaddr_t0 (\tmp_icache_dreq_if_cache.vaddr_t0 ),
  //  .\icache_dreq_o.vaddr_t1 (\tmp_icache_dreq_if_cache.vaddr_t1 ),
  //  .pc_commit_i(pc_commit),
  //  .pc_commit_i_t0(pc_commit_t0),
  //  .pc_commit_i_t1(pc_commit_t1),
  //  .\resolved_branch_i.cf_type (\resolved_branch.cf_type ),
  //  .\resolved_branch_i.cf_type_t0 (\resolved_branch.cf_type_t0 ),
  //  .\resolved_branch_i.cf_type_t1 (\resolved_branch.cf_type_t1 ),
  //  .\resolved_branch_i.is_mispredict (\resolved_branch.is_mispredict ),
  //  .\resolved_branch_i.is_mispredict_t0 (\resolved_branch.is_mispredict_t0 ),
  //  .\resolved_branch_i.is_mispredict_t1 (\resolved_branch.is_mispredict_t1 ),
  //  .\resolved_branch_i.is_taken (\resolved_branch.is_taken ),
  //  .\resolved_branch_i.is_taken_t0 (\resolved_branch.is_taken_t0 ),
  //  .\resolved_branch_i.is_taken_t1 (\resolved_branch.is_taken_t1 ),
  //  .\resolved_branch_i.pc (\resolved_branch.pc ),
  //  .\resolved_branch_i.pc_t0 (\resolved_branch.pc_t0 ),
  //  .\resolved_branch_i.pc_t1 (\resolved_branch.pc_t1 ),
  //  .\resolved_branch_i.target_address (\resolved_branch.target_address ),
  //  .\resolved_branch_i.target_address_t0 (\resolved_branch.target_address_t0 ),
  //  .\resolved_branch_i.target_address_t1 (\resolved_branch.target_address_t1 ),
  //  .\resolved_branch_i.valid (\resolved_branch.valid ),
  //  .\resolved_branch_i.valid_t0 (\resolved_branch.valid_t0 ),
  //  .\resolved_branch_i.valid_t1 (\resolved_branch.valid_t1 ),
  //  .rst_ni(rst_ni),
  //  .set_debug_pc_i(set_debug_pc),
  //  .set_debug_pc_i_t0(set_debug_pc_t0),
  //  .set_debug_pc_i_t1(set_debug_pc_t1),
  //  .set_pc_commit_i(set_pc_ctrl_pcgen),
  //  .set_pc_commit_i_t0(set_pc_ctrl_pcgen_t0),
  //  .set_pc_commit_i_t1(set_pc_ctrl_pcgen_t1),
  //  .trap_vector_base_i(trap_vector_base_commit_pcgen),
  //  .trap_vector_base_i_t0(trap_vector_base_commit_pcgen_t0),
  //  .trap_vector_base_i_t1(trap_vector_base_commit_pcgen_t1)
  //);
  id_stage id_stage_i (
    .clk_i(clk_i),
    .debug_mode_i(debug_mode),
    .debug_mode_i_t0(debug_mode_t0),
    .debug_mode_i_t1(debug_mode_t1),
    .debug_req_i(debug_req_i),
    .debug_req_i_t0(debug_req_i_t0),
    .debug_req_i_t1(debug_req_i_t1),
    .\fetch_entry_i.address (\fetch_entry_if_id.address ),
    .\fetch_entry_i.address_t0 (\fetch_entry_if_id.address_t0 ),
    .\fetch_entry_i.address_t1 (\fetch_entry_if_id.address_t1 ),
    .\fetch_entry_i.branch_predict.cf (\fetch_entry_if_id.branch_predict.cf ),
    .\fetch_entry_i.branch_predict.cf_t0 (\fetch_entry_if_id.branch_predict.cf_t0 ),
    .\fetch_entry_i.branch_predict.cf_t1 (\fetch_entry_if_id.branch_predict.cf_t1 ),
    .\fetch_entry_i.branch_predict.predict_address (\fetch_entry_if_id.branch_predict.predict_address ),
    .\fetch_entry_i.branch_predict.predict_address_t0 (\fetch_entry_if_id.branch_predict.predict_address_t0 ),
    .\fetch_entry_i.branch_predict.predict_address_t1 (\fetch_entry_if_id.branch_predict.predict_address_t1 ),
    .\fetch_entry_i.ex.cause (\fetch_entry_if_id.ex.cause ),
    .\fetch_entry_i.ex.cause_t0 (\fetch_entry_if_id.ex.cause_t0 ),
    .\fetch_entry_i.ex.cause_t1 (\fetch_entry_if_id.ex.cause_t1 ),
    .\fetch_entry_i.ex.tval (\fetch_entry_if_id.ex.tval ),
    .\fetch_entry_i.ex.tval_t0 (\fetch_entry_if_id.ex.tval_t0 ),
    .\fetch_entry_i.ex.tval_t1 (\fetch_entry_if_id.ex.tval_t1 ),
    .\fetch_entry_i.ex.valid (\fetch_entry_if_id.ex.valid ),
    .\fetch_entry_i.ex.valid_t0 (\fetch_entry_if_id.ex.valid_t0 ),
    .\fetch_entry_i.ex.valid_t1 (\fetch_entry_if_id.ex.valid_t1 ),
    .\fetch_entry_i.instruction (\fetch_entry_if_id.instruction ),
    .\fetch_entry_i.instruction_t0 (\fetch_entry_if_id.instruction_t0 ),
    .\fetch_entry_i.instruction_t1 (\fetch_entry_if_id.instruction_t1 ),
    .fetch_entry_ready_o(fetch_ready_id_if),
    .fetch_entry_ready_o_t0(fetch_ready_id_if_t0),
    .fetch_entry_ready_o_t1(fetch_ready_id_if_t1),
    .fetch_entry_valid_i(fetch_valid_if_id),
    .fetch_entry_valid_i_t0(fetch_valid_if_id_t0),
    .fetch_entry_valid_i_t1(fetch_valid_if_id_t1),
    .flush_i(flush_ctrl_if),
    .flush_i_t0(flush_ctrl_if_t0),
    .flush_i_t1(flush_ctrl_if_t1),
    .frm_i(frm_csr_id_issue_ex),
    .frm_i_t0(frm_csr_id_issue_ex_t0),
    .frm_i_t1(frm_csr_id_issue_ex_t1),
    .fs_i(fs),
    .fs_i_t0(fs_t0),
    .fs_i_t1(fs_t1),
    .\irq_ctrl_i.global_enable (\irq_ctrl_csr_id.global_enable ),
    .\irq_ctrl_i.global_enable_t0 (\irq_ctrl_csr_id.global_enable_t0 ),
    .\irq_ctrl_i.global_enable_t1 (\irq_ctrl_csr_id.global_enable_t1 ),
    .\irq_ctrl_i.mideleg (\irq_ctrl_csr_id.mideleg ),
    .\irq_ctrl_i.mideleg_t0 (\irq_ctrl_csr_id.mideleg_t0 ),
    .\irq_ctrl_i.mideleg_t1 (\irq_ctrl_csr_id.mideleg_t1 ),
    .\irq_ctrl_i.mie (\irq_ctrl_csr_id.mie ),
    .\irq_ctrl_i.mie_t0 (\irq_ctrl_csr_id.mie_t0 ),
    .\irq_ctrl_i.mie_t1 (\irq_ctrl_csr_id.mie_t1 ),
    .\irq_ctrl_i.mip (\irq_ctrl_csr_id.mip ),
    .\irq_ctrl_i.mip_t0 (\irq_ctrl_csr_id.mip_t0 ),
    .\irq_ctrl_i.mip_t1 (\irq_ctrl_csr_id.mip_t1 ),
    .\irq_ctrl_i.sie (\irq_ctrl_csr_id.sie ),
    .\irq_ctrl_i.sie_t0 (\irq_ctrl_csr_id.sie_t0 ),
    .\irq_ctrl_i.sie_t1 (\irq_ctrl_csr_id.sie_t1 ),
    .irq_i(2'h0),
    .irq_i_t0(2'h0),
    .irq_i_t1(2'h0),
    .is_ctrl_flow_o(is_ctrl_fow_id_issue),
    .is_ctrl_flow_o_t0(is_ctrl_fow_id_issue_t0),
    .is_ctrl_flow_o_t1(is_ctrl_fow_id_issue_t1),
    .\issue_entry_o.bp.cf (\issue_entry_id_issue.bp.cf ),
    .\issue_entry_o.bp.cf_t0 (\issue_entry_id_issue.bp.cf_t0 ),
    .\issue_entry_o.bp.cf_t1 (\issue_entry_id_issue.bp.cf_t1 ),
    .\issue_entry_o.bp.predict_address (\issue_entry_id_issue.bp.predict_address ),
    .\issue_entry_o.bp.predict_address_t0 (\issue_entry_id_issue.bp.predict_address_t0 ),
    .\issue_entry_o.bp.predict_address_t1 (\issue_entry_id_issue.bp.predict_address_t1 ),
    .\issue_entry_o.ex.cause (\issue_entry_id_issue.ex.cause ),
    .\issue_entry_o.ex.cause_t0 (\issue_entry_id_issue.ex.cause_t0 ),
    .\issue_entry_o.ex.cause_t1 (\issue_entry_id_issue.ex.cause_t1 ),
    .\issue_entry_o.ex.tval (\issue_entry_id_issue.ex.tval ),
    .\issue_entry_o.ex.tval_t0 (\issue_entry_id_issue.ex.tval_t0 ),
    .\issue_entry_o.ex.tval_t1 (\issue_entry_id_issue.ex.tval_t1 ),
    .\issue_entry_o.ex.valid (\issue_entry_id_issue.ex.valid ),
    .\issue_entry_o.ex.valid_t0 (\issue_entry_id_issue.ex.valid_t0 ),
    .\issue_entry_o.ex.valid_t1 (\issue_entry_id_issue.ex.valid_t1 ),
    .\issue_entry_o.fu (\issue_entry_id_issue.fu ),
    .\issue_entry_o.fu_t0 (\issue_entry_id_issue.fu_t0 ),
    .\issue_entry_o.fu_t1 (\issue_entry_id_issue.fu_t1 ),
    .\issue_entry_o.is_compressed (\issue_entry_id_issue.is_compressed ),
    .\issue_entry_o.is_compressed_t0 (\issue_entry_id_issue.is_compressed_t0 ),
    .\issue_entry_o.is_compressed_t1 (\issue_entry_id_issue.is_compressed_t1 ),
    .\issue_entry_o.op (\issue_entry_id_issue.op ),
    .\issue_entry_o.op_t0 (\issue_entry_id_issue.op_t0 ),
    .\issue_entry_o.op_t1 (\issue_entry_id_issue.op_t1 ),
    .\issue_entry_o.pc (\issue_entry_id_issue.pc ),
    .\issue_entry_o.pc_t0 (\issue_entry_id_issue.pc_t0 ),
    .\issue_entry_o.pc_t1 (\issue_entry_id_issue.pc_t1 ),
    .\issue_entry_o.rd (\issue_entry_id_issue.rd ),
    .\issue_entry_o.rd_t0 (\issue_entry_id_issue.rd_t0 ),
    .\issue_entry_o.rd_t1 (\issue_entry_id_issue.rd_t1 ),
    .\issue_entry_o.result (\issue_entry_id_issue.result ),
    .\issue_entry_o.result_t0 (\issue_entry_id_issue.result_t0 ),
    .\issue_entry_o.result_t1 (\issue_entry_id_issue.result_t1 ),
    .\issue_entry_o.rs1 (\issue_entry_id_issue.rs1 ),
    .\issue_entry_o.rs1_t0 (\issue_entry_id_issue.rs1_t0 ),
    .\issue_entry_o.rs1_t1 (\issue_entry_id_issue.rs1_t1 ),
    .\issue_entry_o.rs2 (\issue_entry_id_issue.rs2 ),
    .\issue_entry_o.rs2_t0 (\issue_entry_id_issue.rs2_t0 ),
    .\issue_entry_o.rs2_t1 (\issue_entry_id_issue.rs2_t1 ),
    .\issue_entry_o.trans_id (\issue_entry_id_issue.trans_id ),
    .\issue_entry_o.trans_id_t0 (\issue_entry_id_issue.trans_id_t0 ),
    .\issue_entry_o.trans_id_t1 (\issue_entry_id_issue.trans_id_t1 ),
    .\issue_entry_o.use_imm (\issue_entry_id_issue.use_imm ),
    .\issue_entry_o.use_imm_t0 (\issue_entry_id_issue.use_imm_t0 ),
    .\issue_entry_o.use_imm_t1 (\issue_entry_id_issue.use_imm_t1 ),
    .\issue_entry_o.use_pc (\issue_entry_id_issue.use_pc ),
    .\issue_entry_o.use_pc_t0 (\issue_entry_id_issue.use_pc_t0 ),
    .\issue_entry_o.use_pc_t1 (\issue_entry_id_issue.use_pc_t1 ),
    .\issue_entry_o.use_zimm (\issue_entry_id_issue.use_zimm ),
    .\issue_entry_o.use_zimm_t0 (\issue_entry_id_issue.use_zimm_t0 ),
    .\issue_entry_o.use_zimm_t1 (\issue_entry_id_issue.use_zimm_t1 ),
    .\issue_entry_o.valid (\issue_entry_id_issue.valid ),
    .\issue_entry_o.valid_t0 (\issue_entry_id_issue.valid_t0 ),
    .\issue_entry_o.valid_t1 (\issue_entry_id_issue.valid_t1 ),
    .issue_entry_valid_o(issue_entry_valid_id_issue),
    .issue_entry_valid_o_t0(issue_entry_valid_id_issue_t0),
    .issue_entry_valid_o_t1(issue_entry_valid_id_issue_t1),
    .issue_instr_ack_i(issue_instr_issue_id),
    .issue_instr_ack_i_t0(issue_instr_issue_id_t0),
    .issue_instr_ack_i_t1(issue_instr_issue_id_t1),
    .priv_lvl_i(priv_lvl),
    .priv_lvl_i_t0(priv_lvl_t0),
    .priv_lvl_i_t1(priv_lvl_t1),
    .rst_ni(rst_ni),
    .tsr_i(tsr_csr_id),
    .tsr_i_t0(tsr_csr_id_t0),
    .tsr_i_t1(tsr_csr_id_t1),
    .tvm_i(tvm_csr_id),
    .tvm_i_t0(tvm_csr_id_t0),
    .tvm_i_t1(tvm_csr_id_t1),
    .tw_i(tw_csr_id),
    .tw_i_t0(tw_csr_id_t0),
    .tw_i_t1(tw_csr_id_t1)
  );
  \issue_stage(NR_ENTRIES=32'b0100,NR_WB_PORTS=32'b0100,NR_COMMIT_PORTS=32'b010)  issue_stage_i (
    .alu_valid_o(alu_valid_id_ex),
    .alu_valid_o_t0(alu_valid_id_ex_t0),
    .alu_valid_o_t1(alu_valid_id_ex_t1),
    .\branch_predict_o.cf (\branch_predict_id_ex.cf ),
    .\branch_predict_o.cf_t0 (\branch_predict_id_ex.cf_t0 ),
    .\branch_predict_o.cf_t1 (\branch_predict_id_ex.cf_t1 ),
    .\branch_predict_o.predict_address (\branch_predict_id_ex.predict_address ),
    .\branch_predict_o.predict_address_t0 (\branch_predict_id_ex.predict_address_t0 ),
    .\branch_predict_o.predict_address_t1 (\branch_predict_id_ex.predict_address_t1 ),
    .branch_valid_o(branch_valid_id_ex),
    .branch_valid_o_t0(branch_valid_id_ex_t0),
    .branch_valid_o_t1(branch_valid_id_ex_t1),
    .clk_i(clk_i),
    .commit_ack_i(commit_ack),
    .commit_ack_i_t0(commit_ack_t0),
    .commit_ack_i_t1(commit_ack_t1),
    .\commit_instr_o[0].bp.cf (\commit_instr_id_commit[0].bp.cf ),
    .\commit_instr_o[0].bp.cf_t0 (\commit_instr_id_commit[0].bp.cf_t0 ),
    .\commit_instr_o[0].bp.cf_t1 (\commit_instr_id_commit[0].bp.cf_t1 ),
    .\commit_instr_o[0].bp.predict_address (\commit_instr_id_commit[0].bp.predict_address ),
    .\commit_instr_o[0].bp.predict_address_t0 (\commit_instr_id_commit[0].bp.predict_address_t0 ),
    .\commit_instr_o[0].bp.predict_address_t1 (\commit_instr_id_commit[0].bp.predict_address_t1 ),
    .\commit_instr_o[0].ex.cause (\commit_instr_id_commit[0].ex.cause ),
    .\commit_instr_o[0].ex.cause_t0 (\commit_instr_id_commit[0].ex.cause_t0 ),
    .\commit_instr_o[0].ex.cause_t1 (\commit_instr_id_commit[0].ex.cause_t1 ),
    .\commit_instr_o[0].ex.tval (\commit_instr_id_commit[0].ex.tval ),
    .\commit_instr_o[0].ex.tval_t0 (\commit_instr_id_commit[0].ex.tval_t0 ),
    .\commit_instr_o[0].ex.tval_t1 (\commit_instr_id_commit[0].ex.tval_t1 ),
    .\commit_instr_o[0].ex.valid (\commit_instr_id_commit[0].ex.valid ),
    .\commit_instr_o[0].ex.valid_t0 (\commit_instr_id_commit[0].ex.valid_t0 ),
    .\commit_instr_o[0].ex.valid_t1 (\commit_instr_id_commit[0].ex.valid_t1 ),
    .\commit_instr_o[0].fu (\commit_instr_id_commit[0].fu ),
    .\commit_instr_o[0].fu_t0 (\commit_instr_id_commit[0].fu_t0 ),
    .\commit_instr_o[0].fu_t1 (\commit_instr_id_commit[0].fu_t1 ),
    .\commit_instr_o[0].is_compressed (\commit_instr_id_commit[0].is_compressed ),
    .\commit_instr_o[0].is_compressed_t0 (\commit_instr_id_commit[0].is_compressed_t0 ),
    .\commit_instr_o[0].is_compressed_t1 (\commit_instr_id_commit[0].is_compressed_t1 ),
    .\commit_instr_o[0].op (\commit_instr_id_commit[0].op ),
    .\commit_instr_o[0].op_t0 (\commit_instr_id_commit[0].op_t0 ),
    .\commit_instr_o[0].op_t1 (\commit_instr_id_commit[0].op_t1 ),
    .\commit_instr_o[0].pc (\commit_instr_id_commit[0].pc ),
    .\commit_instr_o[0].pc_t0 (\commit_instr_id_commit[0].pc_t0 ),
    .\commit_instr_o[0].pc_t1 (\commit_instr_id_commit[0].pc_t1 ),
    .\commit_instr_o[0].rd (\commit_instr_id_commit[0].rd ),
    .\commit_instr_o[0].rd_t0 (\commit_instr_id_commit[0].rd_t0 ),
    .\commit_instr_o[0].rd_t1 (\commit_instr_id_commit[0].rd_t1 ),
    .\commit_instr_o[0].result (\commit_instr_id_commit[0].result ),
    .\commit_instr_o[0].result_t0 (\commit_instr_id_commit[0].result_t0 ),
    .\commit_instr_o[0].result_t1 (\commit_instr_id_commit[0].result_t1 ),
    .\commit_instr_o[0].rs1 (\commit_instr_id_commit[0].rs1 ),
    .\commit_instr_o[0].rs1_t0 (\commit_instr_id_commit[0].rs1_t0 ),
    .\commit_instr_o[0].rs1_t1 (\commit_instr_id_commit[0].rs1_t1 ),
    .\commit_instr_o[0].rs2 (\commit_instr_id_commit[0].rs2 ),
    .\commit_instr_o[0].rs2_t0 (\commit_instr_id_commit[0].rs2_t0 ),
    .\commit_instr_o[0].rs2_t1 (\commit_instr_id_commit[0].rs2_t1 ),
    .\commit_instr_o[0].trans_id (\commit_instr_id_commit[0].trans_id ),
    .\commit_instr_o[0].trans_id_t0 (\commit_instr_id_commit[0].trans_id_t0 ),
    .\commit_instr_o[0].trans_id_t1 (\commit_instr_id_commit[0].trans_id_t1 ),
    .\commit_instr_o[0].use_imm (\commit_instr_id_commit[0].use_imm ),
    .\commit_instr_o[0].use_imm_t0 (\commit_instr_id_commit[0].use_imm_t0 ),
    .\commit_instr_o[0].use_imm_t1 (\commit_instr_id_commit[0].use_imm_t1 ),
    .\commit_instr_o[0].use_pc (\commit_instr_id_commit[0].use_pc ),
    .\commit_instr_o[0].use_pc_t0 (\commit_instr_id_commit[0].use_pc_t0 ),
    .\commit_instr_o[0].use_pc_t1 (\commit_instr_id_commit[0].use_pc_t1 ),
    .\commit_instr_o[0].use_zimm (\commit_instr_id_commit[0].use_zimm ),
    .\commit_instr_o[0].use_zimm_t0 (\commit_instr_id_commit[0].use_zimm_t0 ),
    .\commit_instr_o[0].use_zimm_t1 (\commit_instr_id_commit[0].use_zimm_t1 ),
    .\commit_instr_o[0].valid (\commit_instr_id_commit[0].valid ),
    .\commit_instr_o[0].valid_t0 (\commit_instr_id_commit[0].valid_t0 ),
    .\commit_instr_o[0].valid_t1 (\commit_instr_id_commit[0].valid_t1 ),
    .\commit_instr_o[1].bp.cf (\commit_instr_id_commit[1].bp.cf ),
    .\commit_instr_o[1].bp.cf_t0 (\commit_instr_id_commit[1].bp.cf_t0 ),
    .\commit_instr_o[1].bp.cf_t1 (\commit_instr_id_commit[1].bp.cf_t1 ),
    .\commit_instr_o[1].bp.predict_address (\commit_instr_id_commit[1].bp.predict_address ),
    .\commit_instr_o[1].bp.predict_address_t0 (\commit_instr_id_commit[1].bp.predict_address_t0 ),
    .\commit_instr_o[1].bp.predict_address_t1 (\commit_instr_id_commit[1].bp.predict_address_t1 ),
    .\commit_instr_o[1].ex.cause (\commit_instr_id_commit[1].ex.cause ),
    .\commit_instr_o[1].ex.cause_t0 (\commit_instr_id_commit[1].ex.cause_t0 ),
    .\commit_instr_o[1].ex.cause_t1 (\commit_instr_id_commit[1].ex.cause_t1 ),
    .\commit_instr_o[1].ex.tval (\commit_instr_id_commit[1].ex.tval ),
    .\commit_instr_o[1].ex.tval_t0 (\commit_instr_id_commit[1].ex.tval_t0 ),
    .\commit_instr_o[1].ex.tval_t1 (\commit_instr_id_commit[1].ex.tval_t1 ),
    .\commit_instr_o[1].ex.valid (\commit_instr_id_commit[1].ex.valid ),
    .\commit_instr_o[1].ex.valid_t0 (\commit_instr_id_commit[1].ex.valid_t0 ),
    .\commit_instr_o[1].ex.valid_t1 (\commit_instr_id_commit[1].ex.valid_t1 ),
    .\commit_instr_o[1].fu (\commit_instr_id_commit[1].fu ),
    .\commit_instr_o[1].fu_t0 (\commit_instr_id_commit[1].fu_t0 ),
    .\commit_instr_o[1].fu_t1 (\commit_instr_id_commit[1].fu_t1 ),
    .\commit_instr_o[1].is_compressed (\commit_instr_id_commit[1].is_compressed ),
    .\commit_instr_o[1].is_compressed_t0 (\commit_instr_id_commit[1].is_compressed_t0 ),
    .\commit_instr_o[1].is_compressed_t1 (\commit_instr_id_commit[1].is_compressed_t1 ),
    .\commit_instr_o[1].op (\commit_instr_id_commit[1].op ),
    .\commit_instr_o[1].op_t0 (\commit_instr_id_commit[1].op_t0 ),
    .\commit_instr_o[1].op_t1 (\commit_instr_id_commit[1].op_t1 ),
    .\commit_instr_o[1].pc (\commit_instr_id_commit[1].pc ),
    .\commit_instr_o[1].pc_t0 (\commit_instr_id_commit[1].pc_t0 ),
    .\commit_instr_o[1].pc_t1 (\commit_instr_id_commit[1].pc_t1 ),
    .\commit_instr_o[1].rd (\commit_instr_id_commit[1].rd ),
    .\commit_instr_o[1].rd_t0 (\commit_instr_id_commit[1].rd_t0 ),
    .\commit_instr_o[1].rd_t1 (\commit_instr_id_commit[1].rd_t1 ),
    .\commit_instr_o[1].result (\commit_instr_id_commit[1].result ),
    .\commit_instr_o[1].result_t0 (\commit_instr_id_commit[1].result_t0 ),
    .\commit_instr_o[1].result_t1 (\commit_instr_id_commit[1].result_t1 ),
    .\commit_instr_o[1].rs1 (\commit_instr_id_commit[1].rs1 ),
    .\commit_instr_o[1].rs1_t0 (\commit_instr_id_commit[1].rs1_t0 ),
    .\commit_instr_o[1].rs1_t1 (\commit_instr_id_commit[1].rs1_t1 ),
    .\commit_instr_o[1].rs2 (\commit_instr_id_commit[1].rs2 ),
    .\commit_instr_o[1].rs2_t0 (\commit_instr_id_commit[1].rs2_t0 ),
    .\commit_instr_o[1].rs2_t1 (\commit_instr_id_commit[1].rs2_t1 ),
    .\commit_instr_o[1].trans_id (\commit_instr_id_commit[1].trans_id ),
    .\commit_instr_o[1].trans_id_t0 (\commit_instr_id_commit[1].trans_id_t0 ),
    .\commit_instr_o[1].trans_id_t1 (\commit_instr_id_commit[1].trans_id_t1 ),
    .\commit_instr_o[1].use_imm (\commit_instr_id_commit[1].use_imm ),
    .\commit_instr_o[1].use_imm_t0 (\commit_instr_id_commit[1].use_imm_t0 ),
    .\commit_instr_o[1].use_imm_t1 (\commit_instr_id_commit[1].use_imm_t1 ),
    .\commit_instr_o[1].use_pc (\commit_instr_id_commit[1].use_pc ),
    .\commit_instr_o[1].use_pc_t0 (\commit_instr_id_commit[1].use_pc_t0 ),
    .\commit_instr_o[1].use_pc_t1 (\commit_instr_id_commit[1].use_pc_t1 ),
    .\commit_instr_o[1].use_zimm (\commit_instr_id_commit[1].use_zimm ),
    .\commit_instr_o[1].use_zimm_t0 (\commit_instr_id_commit[1].use_zimm_t0 ),
    .\commit_instr_o[1].use_zimm_t1 (\commit_instr_id_commit[1].use_zimm_t1 ),
    .\commit_instr_o[1].valid (\commit_instr_id_commit[1].valid ),
    .\commit_instr_o[1].valid_t0 (\commit_instr_id_commit[1].valid_t0 ),
    .\commit_instr_o[1].valid_t1 (\commit_instr_id_commit[1].valid_t1 ),
    .csr_valid_o(csr_valid_id_ex),
    .csr_valid_o_t0(csr_valid_id_ex_t0),
    .csr_valid_o_t1(csr_valid_id_ex_t1),
    .decoded_instr_ack_o(issue_instr_issue_id),
    .decoded_instr_ack_o_t0(issue_instr_issue_id_t0),
    .decoded_instr_ack_o_t1(issue_instr_issue_id_t1),
    .\decoded_instr_i.bp.cf (\issue_entry_id_issue.bp.cf ),
    .\decoded_instr_i.bp.cf_t0 (\issue_entry_id_issue.bp.cf_t0 ),
    .\decoded_instr_i.bp.cf_t1 (\issue_entry_id_issue.bp.cf_t1 ),
    .\decoded_instr_i.bp.predict_address (\issue_entry_id_issue.bp.predict_address ),
    .\decoded_instr_i.bp.predict_address_t0 (\issue_entry_id_issue.bp.predict_address_t0 ),
    .\decoded_instr_i.bp.predict_address_t1 (\issue_entry_id_issue.bp.predict_address_t1 ),
    .\decoded_instr_i.ex.cause (\issue_entry_id_issue.ex.cause ),
    .\decoded_instr_i.ex.cause_t0 (\issue_entry_id_issue.ex.cause_t0 ),
    .\decoded_instr_i.ex.cause_t1 (\issue_entry_id_issue.ex.cause_t1 ),
    .\decoded_instr_i.ex.tval (\issue_entry_id_issue.ex.tval ),
    .\decoded_instr_i.ex.tval_t0 (\issue_entry_id_issue.ex.tval_t0 ),
    .\decoded_instr_i.ex.tval_t1 (\issue_entry_id_issue.ex.tval_t1 ),
    .\decoded_instr_i.ex.valid (\issue_entry_id_issue.ex.valid ),
    .\decoded_instr_i.ex.valid_t0 (\issue_entry_id_issue.ex.valid_t0 ),
    .\decoded_instr_i.ex.valid_t1 (\issue_entry_id_issue.ex.valid_t1 ),
    .\decoded_instr_i.fu (\issue_entry_id_issue.fu ),
    .\decoded_instr_i.fu_t0 (\issue_entry_id_issue.fu_t0 ),
    .\decoded_instr_i.fu_t1 (\issue_entry_id_issue.fu_t1 ),
    .\decoded_instr_i.is_compressed (\issue_entry_id_issue.is_compressed ),
    .\decoded_instr_i.is_compressed_t0 (\issue_entry_id_issue.is_compressed_t0 ),
    .\decoded_instr_i.is_compressed_t1 (\issue_entry_id_issue.is_compressed_t1 ),
    .\decoded_instr_i.op (\issue_entry_id_issue.op ),
    .\decoded_instr_i.op_t0 (\issue_entry_id_issue.op_t0 ),
    .\decoded_instr_i.op_t1 (\issue_entry_id_issue.op_t1 ),
    .\decoded_instr_i.pc (\issue_entry_id_issue.pc ),
    .\decoded_instr_i.pc_t0 (\issue_entry_id_issue.pc_t0 ),
    .\decoded_instr_i.pc_t1 (\issue_entry_id_issue.pc_t1 ),
    .\decoded_instr_i.rd (\issue_entry_id_issue.rd ),
    .\decoded_instr_i.rd_t0 (\issue_entry_id_issue.rd_t0 ),
    .\decoded_instr_i.rd_t1 (\issue_entry_id_issue.rd_t1 ),
    .\decoded_instr_i.result (\issue_entry_id_issue.result ),
    .\decoded_instr_i.result_t0 (\issue_entry_id_issue.result_t0 ),
    .\decoded_instr_i.result_t1 (\issue_entry_id_issue.result_t1 ),
    .\decoded_instr_i.rs1 (\issue_entry_id_issue.rs1 ),
    .\decoded_instr_i.rs1_t0 (\issue_entry_id_issue.rs1_t0 ),
    .\decoded_instr_i.rs1_t1 (\issue_entry_id_issue.rs1_t1 ),
    .\decoded_instr_i.rs2 (\issue_entry_id_issue.rs2 ),
    .\decoded_instr_i.rs2_t0 (\issue_entry_id_issue.rs2_t0 ),
    .\decoded_instr_i.rs2_t1 (\issue_entry_id_issue.rs2_t1 ),
    .\decoded_instr_i.trans_id (\issue_entry_id_issue.trans_id ),
    .\decoded_instr_i.trans_id_t0 (\issue_entry_id_issue.trans_id_t0 ),
    .\decoded_instr_i.trans_id_t1 (\issue_entry_id_issue.trans_id_t1 ),
    .\decoded_instr_i.use_imm (\issue_entry_id_issue.use_imm ),
    .\decoded_instr_i.use_imm_t0 (\issue_entry_id_issue.use_imm_t0 ),
    .\decoded_instr_i.use_imm_t1 (\issue_entry_id_issue.use_imm_t1 ),
    .\decoded_instr_i.use_pc (\issue_entry_id_issue.use_pc ),
    .\decoded_instr_i.use_pc_t0 (\issue_entry_id_issue.use_pc_t0 ),
    .\decoded_instr_i.use_pc_t1 (\issue_entry_id_issue.use_pc_t1 ),
    .\decoded_instr_i.use_zimm (\issue_entry_id_issue.use_zimm ),
    .\decoded_instr_i.use_zimm_t0 (\issue_entry_id_issue.use_zimm_t0 ),
    .\decoded_instr_i.use_zimm_t1 (\issue_entry_id_issue.use_zimm_t1 ),
    .\decoded_instr_i.valid (\issue_entry_id_issue.valid ),
    .\decoded_instr_i.valid_t0 (\issue_entry_id_issue.valid_t0 ),
    .\decoded_instr_i.valid_t1 (\issue_entry_id_issue.valid_t1 ),
    .decoded_instr_valid_i(issue_entry_valid_id_issue),
    .decoded_instr_valid_i_t0(issue_entry_valid_id_issue_t0),
    .decoded_instr_valid_i_t1(issue_entry_valid_id_issue_t1),
    .\ex_ex_i[0].cause (\fpu_exception_ex_id.cause ),
    .\ex_ex_i[0].cause_t0 (\fpu_exception_ex_id.cause_t0 ),
    .\ex_ex_i[0].cause_t1 (\fpu_exception_ex_id.cause_t1 ),
    .\ex_ex_i[0].tval (\fpu_exception_ex_id.tval ),
    .\ex_ex_i[0].tval_t0 (\fpu_exception_ex_id.tval_t0 ),
    .\ex_ex_i[0].tval_t1 (\fpu_exception_ex_id.tval_t1 ),
    .\ex_ex_i[0].valid (\fpu_exception_ex_id.valid ),
    .\ex_ex_i[0].valid_t0 (\fpu_exception_ex_id.valid_t0 ),
    .\ex_ex_i[0].valid_t1 (\fpu_exception_ex_id.valid_t1 ),
    .\ex_ex_i[1].cause (\store_exception_ex_id.cause ),
    .\ex_ex_i[1].cause_t0 (\store_exception_ex_id.cause_t0 ),
    .\ex_ex_i[1].cause_t1 (\store_exception_ex_id.cause_t1 ),
    .\ex_ex_i[1].tval (\store_exception_ex_id.tval ),
    .\ex_ex_i[1].tval_t0 (\store_exception_ex_id.tval_t0 ),
    .\ex_ex_i[1].tval_t1 (\store_exception_ex_id.tval_t1 ),
    .\ex_ex_i[1].valid (\store_exception_ex_id.valid ),
    .\ex_ex_i[1].valid_t0 (\store_exception_ex_id.valid_t0 ),
    .\ex_ex_i[1].valid_t1 (\store_exception_ex_id.valid_t1 ),
    .\ex_ex_i[2].cause (\load_exception_ex_id.cause ),
    .\ex_ex_i[2].cause_t0 (\load_exception_ex_id.cause_t0 ),
    .\ex_ex_i[2].cause_t1 (\load_exception_ex_id.cause_t1 ),
    .\ex_ex_i[2].tval (\load_exception_ex_id.tval ),
    .\ex_ex_i[2].tval_t0 (\load_exception_ex_id.tval_t0 ),
    .\ex_ex_i[2].tval_t1 (\load_exception_ex_id.tval_t1 ),
    .\ex_ex_i[2].valid (\load_exception_ex_id.valid ),
    .\ex_ex_i[2].valid_t0 (\load_exception_ex_id.valid_t0 ),
    .\ex_ex_i[2].valid_t1 (\load_exception_ex_id.valid_t1 ),
    .\ex_ex_i[3].cause (\flu_exception_ex_id.cause ),
    .\ex_ex_i[3].cause_t0 (\flu_exception_ex_id.cause_t0 ),
    .\ex_ex_i[3].cause_t1 (\flu_exception_ex_id.cause_t1 ),
    .\ex_ex_i[3].tval (\flu_exception_ex_id.tval ),
    .\ex_ex_i[3].tval_t0 (\flu_exception_ex_id.tval_t0 ),
    .\ex_ex_i[3].tval_t1 (\flu_exception_ex_id.tval_t1 ),
    .\ex_ex_i[3].valid (\flu_exception_ex_id.valid ),
    .\ex_ex_i[3].valid_t0 (\flu_exception_ex_id.valid_t0 ),
    .\ex_ex_i[3].valid_t1 (\flu_exception_ex_id.valid_t1 ),
    .flu_ready_i(flu_ready_ex_id),
    .flu_ready_i_t0(flu_ready_ex_id_t0),
    .flu_ready_i_t1(flu_ready_ex_id_t1),
    .flush_i(flush_ctrl_id),
    .flush_i_t0(flush_ctrl_id_t0),
    .flush_i_t1(flush_ctrl_id_t1),
    .flush_unissued_instr_i(flush_unissued_instr_ctrl_id),
    .flush_unissued_instr_i_t0(flush_unissued_instr_ctrl_id_t0),
    .flush_unissued_instr_i_t1(flush_unissued_instr_ctrl_id_t1),
    .fpu_fmt_o(fpu_fmt_id_ex),
    .fpu_fmt_o_t0(fpu_fmt_id_ex_t0),
    .fpu_fmt_o_t1(fpu_fmt_id_ex_t1),
    .fpu_ready_i(fpu_ready_ex_id),
    .fpu_ready_i_t0(fpu_ready_ex_id_t0),
    .fpu_ready_i_t1(fpu_ready_ex_id_t1),
    .fpu_rm_o(fpu_rm_id_ex),
    .fpu_rm_o_t0(fpu_rm_id_ex_t0),
    .fpu_rm_o_t1(fpu_rm_id_ex_t1),
    .fpu_valid_o(fpu_valid_id_ex),
    .fpu_valid_o_t0(fpu_valid_id_ex_t0),
    .fpu_valid_o_t1(fpu_valid_id_ex_t1),
    .\fu_data_o.fu (\fu_data_id_ex.fu ),
    .\fu_data_o.fu_t0 (\fu_data_id_ex.fu_t0 ),
    .\fu_data_o.fu_t1 (\fu_data_id_ex.fu_t1 ),
    .\fu_data_o.imm (\fu_data_id_ex.imm ),
    .\fu_data_o.imm_t0 (\fu_data_id_ex.imm_t0 ),
    .\fu_data_o.imm_t1 (\fu_data_id_ex.imm_t1 ),
    .\fu_data_o.operand_a (\fu_data_id_ex.operand_a ),
    .\fu_data_o.operand_a_t0 (\fu_data_id_ex.operand_a_t0 ),
    .\fu_data_o.operand_a_t1 (\fu_data_id_ex.operand_a_t1 ),
    .\fu_data_o.operand_b (\fu_data_id_ex.operand_b ),
    .\fu_data_o.operand_b_t0 (\fu_data_id_ex.operand_b_t0 ),
    .\fu_data_o.operand_b_t1 (\fu_data_id_ex.operand_b_t1 ),
    .\fu_data_o.operator (\fu_data_id_ex.operator ),
    .\fu_data_o.operator_t0 (\fu_data_id_ex.operator_t0 ),
    .\fu_data_o.operator_t1 (\fu_data_id_ex.operator_t1 ),
    .\fu_data_o.trans_id (\fu_data_id_ex.trans_id ),
    .\fu_data_o.trans_id_t0 (\fu_data_id_ex.trans_id_t0 ),
    .\fu_data_o.trans_id_t1 (\fu_data_id_ex.trans_id_t1 ),
    .is_compressed_instr_o(is_compressed_instr_id_ex),
    .is_compressed_instr_o_t0(is_compressed_instr_id_ex_t0),
    .is_compressed_instr_o_t1(is_compressed_instr_id_ex_t1),
    .is_ctrl_flow_i(is_ctrl_fow_id_issue),
    .is_ctrl_flow_i_t0(is_ctrl_fow_id_issue_t0),
    .is_ctrl_flow_i_t1(is_ctrl_fow_id_issue_t1),
    .lsu_ready_i(lsu_ready_ex_id),
    .lsu_ready_i_t0(lsu_ready_ex_id_t0),
    .lsu_ready_i_t1(lsu_ready_ex_id_t1),
    .lsu_valid_o(lsu_valid_id_ex),
    .lsu_valid_o_t0(lsu_valid_id_ex_t0),
    .lsu_valid_o_t1(lsu_valid_id_ex_t1),
    .mult_valid_o(mult_valid_id_ex),
    .mult_valid_o_t0(mult_valid_id_ex_t0),
    .mult_valid_o_t1(mult_valid_id_ex_t1),
    .pc_o(pc_id_ex),
    .pc_o_t0(pc_id_ex_t0),
    .pc_o_t1(pc_id_ex_t1),
    .resolve_branch_i(resolve_branch_ex_id),
    .resolve_branch_i_t0(resolve_branch_ex_id_t0),
    .resolve_branch_i_t1(resolve_branch_ex_id_t1),
    .\resolved_branch_i.cf_type (\resolved_branch.cf_type ),
    .\resolved_branch_i.cf_type_t0 (\resolved_branch.cf_type_t0 ),
    .\resolved_branch_i.cf_type_t1 (\resolved_branch.cf_type_t1 ),
    .\resolved_branch_i.is_mispredict (\resolved_branch.is_mispredict ),
    .\resolved_branch_i.is_mispredict_t0 (\resolved_branch.is_mispredict_t0 ),
    .\resolved_branch_i.is_mispredict_t1 (\resolved_branch.is_mispredict_t1 ),
    .\resolved_branch_i.is_taken (\resolved_branch.is_taken ),
    .\resolved_branch_i.is_taken_t0 (\resolved_branch.is_taken_t0 ),
    .\resolved_branch_i.is_taken_t1 (\resolved_branch.is_taken_t1 ),
    .\resolved_branch_i.pc (\resolved_branch.pc ),
    .\resolved_branch_i.pc_t0 (\resolved_branch.pc_t0 ),
    .\resolved_branch_i.pc_t1 (\resolved_branch.pc_t1 ),
    .\resolved_branch_i.target_address (\resolved_branch.target_address ),
    .\resolved_branch_i.target_address_t0 (\resolved_branch.target_address_t0 ),
    .\resolved_branch_i.target_address_t1 (\resolved_branch.target_address_t1 ),
    .\resolved_branch_i.valid (\resolved_branch.valid ),
    .\resolved_branch_i.valid_t0 (\resolved_branch.valid_t0 ),
    .\resolved_branch_i.valid_t1 (\resolved_branch.valid_t1 ),
    .rs1_forwarding_o(rs1_forwarding_id_ex),
    .rs1_forwarding_o_t0(rs1_forwarding_id_ex_t0),
    .rs1_forwarding_o_t1(rs1_forwarding_id_ex_t1),
    .rs2_forwarding_o(rs2_forwarding_id_ex),
    .rs2_forwarding_o_t0(rs2_forwarding_id_ex_t0),
    .rs2_forwarding_o_t1(rs2_forwarding_id_ex_t1),
    .rst_ni(rst_ni),
    .sb_full_o(sb_full),
    .sb_full_o_t0(sb_full_t0),
    .sb_full_o_t1(sb_full_t1),
    .\trans_id_i[0] (fpu_trans_id_ex_id),
    .\trans_id_i[0]_t0 (fpu_trans_id_ex_id_t0),
    .\trans_id_i[0]_t1 (fpu_trans_id_ex_id_t1),
    .\trans_id_i[1] (store_trans_id_ex_id),
    .\trans_id_i[1]_t0 (store_trans_id_ex_id_t0),
    .\trans_id_i[1]_t1 (store_trans_id_ex_id_t1),
    .\trans_id_i[2] (load_trans_id_ex_id),
    .\trans_id_i[2]_t0 (load_trans_id_ex_id_t0),
    .\trans_id_i[2]_t1 (load_trans_id_ex_id_t1),
    .\trans_id_i[3] (flu_trans_id_ex_id),
    .\trans_id_i[3]_t0 (flu_trans_id_ex_id_t0),
    .\trans_id_i[3]_t1 (flu_trans_id_ex_id_t1),
    .\waddr_i[0] (\waddr_commit_id[0] ),
    .\waddr_i[0]_t0 (\waddr_commit_id[0]_t0 ),
    .\waddr_i[0]_t1 (\waddr_commit_id[0]_t1 ),
    .\waddr_i[1] (\waddr_commit_id[1] ),
    .\waddr_i[1]_t0 (\waddr_commit_id[1]_t0 ),
    .\waddr_i[1]_t1 (\waddr_commit_id[1]_t1 ),
    .\wbdata_i[0] (fpu_result_ex_id),
    .\wbdata_i[0]_t0 (fpu_result_ex_id_t0),
    .\wbdata_i[0]_t1 (fpu_result_ex_id_t1),
    .\wbdata_i[1] (store_result_ex_id),
    .\wbdata_i[1]_t0 (store_result_ex_id_t0),
    .\wbdata_i[1]_t1 (store_result_ex_id_t1),
    .\wbdata_i[2] (load_result_ex_id),
    .\wbdata_i[2]_t0 (load_result_ex_id_t0),
    .\wbdata_i[2]_t1 (load_result_ex_id_t1),
    .\wbdata_i[3] (flu_result_ex_id),
    .\wbdata_i[3]_t0 (flu_result_ex_id_t0),
    .\wbdata_i[3]_t1 (flu_result_ex_id_t1),
    .\wdata_i[0] (\wdata_commit_id[0] ),
    .\wdata_i[0]_t0 (\wdata_commit_id[0]_t0 ),
    .\wdata_i[0]_t1 (\wdata_commit_id[0]_t1 ),
    .\wdata_i[1] (\wdata_commit_id[1] ),
    .\wdata_i[1]_t0 (\wdata_commit_id[1]_t0 ),
    .\wdata_i[1]_t1 (\wdata_commit_id[1]_t1 ),
    .we_fpr_i(we_fpr_commit_id),
    .we_fpr_i_t0(we_fpr_commit_id_t0),
    .we_fpr_i_t1(we_fpr_commit_id_t1),
    .we_gpr_i(we_gpr_commit_id),
    .we_gpr_i_t0(we_gpr_commit_id_t0),
    .we_gpr_i_t1(we_gpr_commit_id_t1),
    .wt_valid_i({ flu_valid_ex_id, load_valid_ex_id, store_valid_ex_id, fpu_valid_ex_id }),
    .wt_valid_i_t0({ flu_valid_ex_id_t0, load_valid_ex_id_t0, store_valid_ex_id_t0, fpu_valid_ex_id_t0 }),
    .wt_valid_i_t1({ flu_valid_ex_id_t1, load_valid_ex_id_t1, store_valid_ex_id_t1, fpu_valid_ex_id_t1 })
  );
  assign _9292_ = 1'h0;
  assign _9295_ = 1'h1;
  assign irq_i = 2'h0;
  assign boot_addr_i = 64'h0000000000000000;
  assign hart_id_i = 64'h0000000000000000;
  assign no_st_pending_commit_t0 = no_st_pending_ex_t0;
  assign no_st_pending_commit_t1 = no_st_pending_ex_t1;
  assign dcache_flush_ack_cache_ctrl_t0 = 1'h0;
  assign dcache_flush_ack_cache_ctrl_t1 = 1'h0;
  assign ipi_i_t0 = 1'h0;
  assign ipi_i_t1 = 1'h0;
  assign time_irq_i_t0 = 1'h0;
  assign time_irq_i_t1 = 1'h0;
  assign debug_req_i_t0 = 1'h0;
  assign debug_req_i_t1 = 1'h0;
  assign _9293_ = 1'h0;
  assign _9294_ = 1'h0;
  assign _9296_ = 1'h0;
  assign _9297_ = 1'h0;
  assign irq_i_t0 = 2'h0;
  assign irq_i_t1 = 2'h0;
  assign boot_addr_i_t0 = 64'h0000000000000000;
  assign boot_addr_i_t1 = 64'h0000000000000000;
  assign hart_id_i_t0 = 64'h0000000000000000;
  assign hart_id_i_t1 = 64'h0000000000000000;
endmodule
