i_SW_0: assume property (i0[14:12] == 3'b010);
i_SW_1: assume property (i0[6:0] == 7'b0100011);
