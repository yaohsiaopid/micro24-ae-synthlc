group_14_i0: assume property (
(i0[31:28] == 4'b0000 && i0[27:24] == 4'b0000 && i0[23:20] == 4'b0000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b001 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b0001111 &&  1'b1 ) || 
(i0[31:28] == 4'b0000 && i0[19:15] == 5'b00000 && i0[14:12] == 3'b000 && i0[11:7] == 5'b00000 && i0[6:0] == 7'b0001111 &&  1'b1 ) || 
1'b0);
//14||FENCE,FENCEI
