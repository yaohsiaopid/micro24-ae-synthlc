`define SYSINSN
i_CSRRCI_0: assume property (i0[14:12] == 3'b111);
i_CSRRCI_2: assume property (i0[6:0] == 7'b1110011);
